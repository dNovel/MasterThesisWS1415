MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���eܻ�eܻ�eܻ+D��eܻ��B��eܻ��v��eܻ�O��eܻ�eݻ�eܻ��w��eܻ��G��eܻ��A��eܻRich�eܻ        PE  L ��P        � !
  n	  �     �                             �                             0 b   ` (                            p LC  `�                                            �a �                          .textbssUk                        �  �.text   Km	  �  n	                   `.rdata  �  �    r	             @  @.data   ,E        �
             @  �.idata  	   `     �
             @  �.reloc  O   p  P   �
             @  B                                                                                                                                                                                                                                                                                                                        ������l �q �� �w� �� �� �>8	 ��� �NW ��� �� 鿷 �z ��f �	 �@ �&2 ��� �� �U � �]� ��� ��� �� ��� �*	 ��H ��  �E	 ��� �{ ��� �!� �l� �. �� �= �� 飭  ��� �ig �	 �D �*	 �y 逽 �Kf ��: �� �� �6 颇 �m� �l7	 �c� �? �Y�  ��o �?�  �z �H ���  �Q �6� �a  ��p ��� ��� �}� �^ �Ө �n� ��Z �T�  �?� �:	 饩 �g ��� ��T �q� �� �7D �{ �]� 騂 ���  �; �� �4y �" ��R �x � � �k$ �v0 �% �\Z �Ǽ  �"j �ݤ �� ��  �޲ �yS �Ե �	 �� �eZ � � �& ��� �Qx ��,	 ��5	 ��� �]� �h�  �� �~` �9�  �Ĭ ��� �Z: �w �p4 ��� �V( ��4 ��# �, �K �} �L ��? ��� �i� �@ �� �K �%�  � �; ��  �aJ 鼡 ��O ��  ��T �(g �C) �N�  �ɫ ��  ��� ��� �գ  �� �۽ � ��� �l	 �g ��N 魍 ��� �c�  �nZ �r �� �� �*  �%m �a �k �Fd �q� �<� �h �M �g  �H�  �j �. �4 �d ���  ��Q �5� �� �+; �f� � �\` ��  �b� 靘 �x� �3l �� ��� ��I �� �J	 ��! �0� �[j 鶻  �ч  �l, �W� �� �=# ��3	 ��� �>f �ɼ ��F �3	 �J� �8 �к  �+ �:5	 � 鼑 �� �b� �-	 �H9 ��6 �.� �)�  �$� �� �� ��� �0$ ��  �6�  �� �\; �� �� ��� �� �3	 ��: �)p 鄙 �� ��� �d �` 黎  �/ �� �T �� 颃 �� 騧 �s� �N� ��� �$ �
 �z� �� �p� ��  ��� �! ��3	 �w< �Ң ��i �� �S	 �; �yv �� ��  �Z� �e  ��  ��L �f �� ��� �� �b� ��� �[ �#W �>� �Y� �A � �Z� �7 ��. 雅  �^ �� �,	 �G1 �R� �m� �/ �c� �>� �� �2	 �O� 隫  �33	 �2 �c �� �# �l# �w � �  �� �S� �>X ��� �T_ �� �3	 酻  �P� � ��� ��a �l, �� �b� ��  � �s 龨 � �t� �=2	 �� �eO �� �[� �f� �Q�  �V �'� �� �� ��� �c/ �n �	� 锔 �O�  �� 饧 �J ��� �6� ��N �L� �� ��M �-
	 鈲 铊 ��  �y~ ��- �� �j� �0	 �`� �[� �F �j� �L. ��� �" ���  騼 �C �� 驱 �j �< 鯬 �e� �@o �+ �v 鑻  �0	 �� 邒 �m� ��� �S �^% �	 ��z �?� �ʵ  �� �` �g1	 ��� �a� �<� �� �K �q ��' ��V ��	 �� ��� ��  �	 饼 ��� �
 ��? ��  ��� �wZ �2� �� �H| �#�  ��� �9� �t� �z �j� ��b ��� �� �ve �� �Lc �W� �B �� �� ���  ��2 �� 鴙 ��� ��� �e� �� �K� �� �� �L� �', �! � �� �
	 �8 �Y1 ���  �_ �� �� � � �{ �V� �� �, �'� �B& �W ��� �3�  �� �9� �� �/� � �ee �� �6 馲  鱦 �|' �g � �J �d.	 � �n� �i� �	 �Ϭ �J�  �%� �0g �� ��-	 �q� ���  ��-	 ��� �m� �X� �3M ��  �	� �� ��a �k 饆 �0� �� �= �A� �� �Ǜ 邴 �� ��= �� ��  �i� ��  � �� �E �S �(	 馫 �a~ 錦 �G� ��u ��� �غ 飩  �Θ  �P ��D �_ 隼 �5� �`X 雜 �&� �!� �L� ��U � �]� �h  铱 �.� ��6 �` �/�  麿 �E� �0� ��  �6�  �; �� �'� �RZ ��� �x� �,	 ��e �Y� �n �?F � �/-	 頇 �[8 �F�  �� �8 �G �� � � ��! �F �% �& ��	 ��� �� 鐈 ��� 閤 �1� �<X �GF �� ��� �X�  �� �h �� �T� ��� �*�  ��� �P ��	 �6� �� �� ��� �� �m 阘 �S � �� ��  ��� 銇 ��� �P�  �+� ��  �A� �,� �G" �� ��  �H� �c� �u �I� �tz �_ �Z�  ���  �p� �k� ��� �A  霴 �g 颱 �X �  �s�  �e �) �- 鏔  �:� �5L �f 鋓 ��h �! �,�  �'# ��� ��� �xv �ӱ �N� ��� �$� ��+	 �� �x �� �[� 醞 �+� 霵 �G� � �s*	 �� �Õ ��O �y�  �2 �_- �
 ��� �� �K �	 ��� �,� �! �� ��� �X� �C� ��y ��% �� 鏆  �H*	 ��6 ��1 ��  �N �1] �|�  �W� � 魫 �� � �.�  ��  �$� ��- ��  �E� ��v �{ �Fw 鱊 �� �g� �rg �� ���  ��*	 �އ  �y2 �� �?� �
� �� �(*	 �+` ��m �
 �, 駧 �R� �� �، �� �W �� ��D �/	 ��� �g �� � ��X � �r*	 �g� �B� 靌 �HC �C� �� �9� �T �O�  �z� �UB �u �k �v� ��  �l �GY �(	 �-b ��� �A 鎙 �Y �dp �/ �:�  �	 �p� 鋔 �
 �� 錂 �)	 �b� �M 阨 �F �^�  ��� �T$ �� �: � �@� �k�  ���  �!� �|� �gs ��P �D �H � �] �� � �/� �Zx �ś �p�  �{� �v� �Ѣ ��y ��` �"� �}Q �� �� �.~ �)s �Ķ  �/� �� �5� ��0 �{� �V� �R ��� ��	 �� �� �H �s� ��� 鹈  �� � �� �& �`� �Ku �f� �� �q ��  �R# ��= 鸸 �s �: �	 �� ��� �:� �� ���  �� �6n  ��u �l	 ��l �� �� �8� �#� �\ ��/ �� �C �:[ �Ÿ �pk �K- �� �ѥ 鼘 �wl  � 	 ��^ �R �� �~ �i� �Դ �Q&	 �*	 �eZ �� �k� �F1 �� �o �� �b	 �� 	 �'	 �3� �� �I/ �T� �� ��� �Ն � � �� �� �, �LS ���  �� �m�  �h�  �C� �_ �1 ��� �C �� ��� ��� �� �� ��9 �� � ���  �]� �H�  �3 �N� ��a �$� �� �z� �U� �� 電  �, �Q} �<� �'� 颰 �-� �� �3; 鎬 �\ �t� 韓  �  ��E ��� �� �ֹ �Q �̣ ��E ��
 �ME �8l ��  �f �)� �t �� 骱 �u ��� ��� ��4 �� ��� �� �"  �M� ��  郔 ��M �* ��� �� �) �u� ��9 髳 �6l � �\� �< � �=� �x! 飪 �Ι � �t �' �ʗ  镯 �P� �;�  �r �� �* ���  �_  ��� �xu ��� �. �i�  �t� ��� �A �� �F �k�  �&e �T �R �w� �2� �B ��� ��Q �� �i� �dp �_� �� �E� � ��o �V�  �� ��� �� �"� �� �L �� �n" ��� � �> � �� � $	 �{� �v� �Q[ �l �' �" �-� �x#	 �C� �� ��r �� ���  ��� �E` �= �� �` �� �  �h �RZ 靑 �h� ��  �N� �� �ԋ �� �� �e� �P �M �& �ё �l� �� �B �ͬ  �8 ��  �~� �i  �� �o �#	 鵂 � � 髞 �fT  �a� �LP �S �
#	 �< �� �L �� �\ �� �O� �ju �5; �z 黨 馢 ��[ � � �` �]� �(# �# �~k �Y� 锛 ���  隽  �� �� �[� �֜ �A{ �"	 �'� �r� � �j �� �ޕ ��! �Ծ �C �J� ��g 逩 鋪 �� �q �,� �v � ��� ��| �C� �( �� �$� �H �
~ � �@Z �[c 閙 �� �!	 釯 ��!	 齼 �h� �CP �v ��) �4j �Ϟ �*g  饓 鰏 �. ��  �� ��8 �G� �br ��t ��� ��� �1 �)� ��  韢 ��  �}!	 鰛 �;A �Fl �1H �� �� �� �e  �4� �#} �>� �9� �t� ���  ��{ �{  �Г �+�  �*!	 �� �� �'� ��  �� ��� ��h ��� �ً �d) ���  �Z8 镾 �0� � �6d � �l� �� �2N �m� �ؾ �#w ��� �y� ��� � �z� �" ��E �[� �v�  �� �<� �� �"� ��� �� �Ü ��� ��� �;� ��� �� �e� �`( �;� �vS �1� �L� 駵 �Ry �� �� �3� �^� 驣  鄔 �? �m  ��/ �PL � �o ��Q ���  ���  �R�  �M� �x� ��c �� �) �- �Q �ڿ �� �p$ �;x ��� �Q�  �<� �� �B" �M �X8 ��( �ޑ �� �dw �3 ��}  ��� �@� 鋿 �
 �	 �� � �� �� �h� �S�  �U �y! � �M �r  ��u  �� �$ �V�  �a�  ��  �W� �"� �� �% �t  �8	 �y( �� �?< 銰 �I �`� ��P ��& �_ �7 ��� �B� �� �g ��d �~? � �� �_ ���  �� �`\ ��� � � �,� �'X �K ��T ��� �� �Ξ �Y0 ��� ��H �*� �e� 鐷 �{k �X  �i	 �� �G� �b  �j �x 铧  �^� �y] �/ �OP �ڒ �5H �p{ �� �&� ��H ��h ���  钷  魊 �p �cS ��  ��� �� �o�  �zy  � ��  �;� �F� �A� �e �� �� � �8 �� �� �	 �$J  �OU ��E � ��� �� �V �1 �<� �w� ��E �� �h	 �� �^y  �X �b  �� ��P  ���  �� �[� ��s �� ��[ �g� �2v �=� �� �2 �nY �) �tL �3 �( �e� � D �  �&y �!� �,� �2 �R? �M� ��? 鳤 ��  �� 锤  �� �jM ��	 �� �+� �vr  ��. �,� �� �� �Q �� 铍 �~] �Y� �� �� �j� ��n � �  ��V �&v ��3 ��  �� �bq �M  ��	 �n 鎘 �Y4 �t: ��  �J� �� � �  �+�  �� �� � �' �� � 鸰 �ӆ ��� �I� �T� � �Z� �� �` ��P �&2 �4 �i �g� �b� �͎ �XE �c� �~� �9 �	 ��  �B �� � ) 黉 � ��� � �  �R� ��e ��  鳼 �^� �9� ���  �_�  �k �U� �`� ��* ��� 遯 �̦ �G� �J 靳 �? �c� �^( �	 �P �M  �Z� �e� ��� 黳 �F ��  �<�  �G� �b\ �Mu ��� �Ct �N� �b ��
 �� �
� �& � �k� �: �4 �4 ���  ��H �͢ �H^ �3, �<	 �9� ��� �� �� �խ �`7 �{s  �V ��{ ��  ��	 �X ��l 鈛 ��I �n �	5 �� �X �:n �?	 鐉 ��F �| 釿 �� ��/ �B� �P �! ��� � ���  �� �  �	 �%� �} ��y �F� �� ��� �h �"� �mY �� �#� �^� �y� �T� �o  ��A �%� �] �} � �� ��! �� �r�  �M� �H �s� 龰 �	� �i� �� �ʴ ��� �@� �;� �? �� �l� ��� �b� �-� � �S� �� �y� �4% �O� ��� � �� �� �� �A�  �� �7� �R
 �m! �� ��- �ާ �Y" �D6 �?� �Z� ��v �� ��� �&� �!� �� ��� �; �]� �� �S� 龯 �W 餾  �_}  �J� �U� �� �� �֊ ��h �\� �w� ���  �� �X� �2 � �9� �S  �� �� �E� �B �k� �f� �!� ��� �G� �� �MU �� �^ 鞒  �i�  �h 鿹 �*� �Z �p� �;� ��M �A�  ��	 �v �b� �� �X8 �S�  ��^ �Y� �� �o� �2 ���  鐰 ��K � �!� �\ �g� �J  ��	 ��� �#G �>h  �� ��\ �/z �� �E� �T	 �� �� �! ��� �
 �R? �� �h �3� �" 际 餵 �O �:�  �Ek  �� ��8 �6� 鑋 �� �� ��I �  �� �#� �n� �
 �d� �� �T	 �%i �I �+� �֋ �q� ��  �y	 �n	 �7 � �#| ��� � �4� �?7 �Zb �ŭ 逭  �{� �v< �Q/ �f �'_ �B@ ��� �Hh  ���  �N7 �I� �D� ��{ �D	 �u�  ��I  �{� �V �k ��5 闎 �b �i  ���  �3I ��� �I� � ��	 ��z �O ��|  ��X  ��� ��� �L� �� 鲋 �}s �h� �3 ��  �� �$� �� 隸 �� �� �� ��  �AO  �� �g# � �-�  �H< �V �Ν �i  �4
 �� �Z� ��  �! �w �fG �� �<) ��� �t  �s 鈧  ��	 �{ � �d�  �� ��� �E	 � � �� ��z ��� �\� �'� �b 靵 �� �#� �q 陲 �� � �
� ��> �0 �+� �&� �� ��� �G� ��/ 齰 ��' �s3 �> �w  �d� ��� 麵 �eg �p		 ��� �&# �� �l � �R 鍄 ��2 �s�  �>� �IC ��� �E �Z� �% ��B  � �v� ��� ��� �x  ��| �: 阴 ���  鎯 ��� �4� ���  �� ��� �P� �+� ��3 �& �R	 ��� �B�  ��J  � �� 鎫 �i) �� �G	 �z� ��C � � �K� �` ��D  �	 釸 ��� �� �8g �C� �n� �� ��� �_�  �� �U� 鐝  �{v ��u �� �	 �W� ��X �] �9 ��k  �L  �z �t � �Q �� ��� �+T �h �� �� ��? �� �-� �h� �� �s �i� �T] ��U 隡  �	 �0� �� � �Q3 ��� ��� �B� ��  ��	 �c� �� �i� �� �� �j� ��  �� ��� �P �a �h	 鷯 � �� �xZ �3� �� �i� �; �_� �& ��  �`�  黸  �fm  �1� �� �W� �B� �݂ ��� �z �~^  �I@ �� �� �� �e� � ���  �6� �aD ��  �e 鲠 �& �v �c� 鮄 ��� ��� �ou 銞  鵵 ��� 髦 �&t �� �$ � �2� ��V �Ȭ  �v 鮻 �	b �4�  � �Z< �E �� �� �� �$ 鼻 �v ��� 鍄 �(� �� �; �r  �� �?� �� �u � L �� 馩 �1 ��h ��� �2� 齂 �5 ��  �^�  ��	 �$� �o� ��: �u{ ��� �� �f� �Q� �( �W� �R� 鍁 �H  �Sa � ��	 ��K �_� �(	 �eq �0� ��� �6# �a
 錫 �wy �b�  �� �� ��� �� ��� �Է �� 銁 �F ��� �[� �6� �	 �� �� �b� �m� �xP ��� �� ��G  �h �?� �*� �UE � � � ��� 顴 �L �L �� �ͫ �� ��� �N� ���  锻  鏯 �*{ �� �@m  �;� �f| �� �P �G� �B� �	 �Ȝ �S �� �Y �$� ��< �Z� ��3 �� ���  ��H ��� �} �G �B� 齾 �h9  �� ��� �Ie �$" �o� �ZL �%� �`�  �� �� �Q� �<L �	 �"Y �e �hi �� �~X �	� �d � �� ��� �`� �� �s �� �,+ �; �2� �� ��	 �s� �� �	j 鄓 �j �:Z  �� �p# �[h �� ��� � ��  题 �}& �X� �S �� �� 齲 �x �*g ��� �F ��� ��� �ѯ �� �s �� ��x �Xl �6 � �� �TI �� �Z�  �u� � Q �[# �� �!� �C  �� �"] ��� �X� �SH �~� 鹦 ��h ��s �:$ �  �`W �a �v ��� �w ��h �� ��� � 
	 �#� ��7  �e �4 �� �
� �ե ��� 髪  �6L �X ��  ���  �n �m�  �� �#� �N� �y	 �tf �_6 �? �1 �0� ���  �� �1� �w  �7 ��f  � �� �� ��� ��  �TH �_� �*� �5�  �F  �u �Vf  ��- �		 �g{ �b~ �=� �x� �� �� �Y�  ��U �� �
 �u� �0� � �	 �� �S �G/ �R 青 阜 �c�  �>� �� �� �S �L		 ��� ��� �� �T �l  �\� ��  �k  �� ��  �1 ��} �Y� �$^ ��H �
 �5� �n  � �F�  �� �,, �$ � � �(� ��� 鎔 �] �4 �_Q  �� 镜  � � �	 醮 �:  ��  ��� �2�  �ݽ �Xy �à �_ ��u �$� ��  �� 饰 ��P �ۜ �ƍ �a� �x � �� �}� ��  ��� �~ �yF �4�  ���  �[ �� �� �[K ��} �< ���  �Y 鲟 �6 �w �� ��� �9	 �D� �� �j� ��� �p� �{� ��  �� �i �W� �¨ �}� ��� �; �N �)� ��u ��  �z� �uu ��� �ۑ ��  ��� �\� �	 �� �-� ��  �	 �~� �	� �]  �_ �z! 饉  � 	 黉 鶣 �q� � �� �o �}� 阹 �3� �N ��t �4c �O! �
� � �p� ��m ��  �� �<� � �2� ��{ �� � �  �	� ��0 ��m �9 ��F �0b  ��  �X  �� ��	 �_ �9 齖 �X�  �� �n�  �	 ��O �?� �9 �� ���  �A 醸 �q� �� �w;  �o �M �X� 郸 �� �9 �t�  �� ��� �^ �P� ���  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E���Ex��M�U;��Զ���EE�E��_^[���   ;�蹶����]� �����������������������U����   SVW��@����0   ������=�* t��EP��*��;��_���_^[���   ;��O�����]��������������������������������U���   SVW��������   ������j h������������P�˟�����E��������c����}� u��  j h��������׿��P�E�P�(�����������������(��������� t�  j h���� ���虿��P�`������E썍 ���������M��՛��j h����P����h���P��8���������8���Pj�M�輷����8���������P�������j h|��������#���P��h����:�����h���Pj�M��w�����h���調���������_���j�������]���������Pj�M��C����������v���j h��������赾��P�������̛��������Pj�M��	����������<���������������}� t1�E�P������蘝���M�Q������Rj�M�趺��������������+�E�P�������g���������Qj�M�蜶���������Ͼ���M������R��P�x�蠟��XZ_^[��   ;�������]�   ������   ��sc �����������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;�������EPj��MQ�U�R��*�H�Q�҃�;��Ĳ���E�_^[���   ;�豲����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;��;���_^[���   ;��+�����]����������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��*���   �H$�у�;��Q����E�_^[���   ;��>�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��*���   �H0�у�;�豰���E�_^[���   ;�螰����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   ��Ѓ�;��)���_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;�贯��_^[���   ;�褯����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M����   ��;��1���_^[���   ;��!�����]� �������������������������������U����   SVW��@����0   �����󫡘*���   ��*��*ǀ�   ͭ蓬����u3���   _^[���   ;�蜮����]�����������������������������U����   SVW��@����0   ������_^[��]������������U���`  SVW�������X   ������E�������������  #�������  tZ������ tB������t�  �������  �u  ��  ��*肔����u3���  �   ��  �   ��  ��  �E�E��E�    �	�E���E�E��M�;�  �E��H�U�<� u��h@��E��H�U��P��������th8��E��H�U��P�Ǜ������u1j h ��������=���������P�\����������������   h��E��H�U��P�x�������u>�E��H�U���    j h ��������޶��������P��������������3����8h���E��H�U��P��������u�E��H�U���    �    �  ������   �E�E��} u�s�E��x t�hj h���������U���������P�M��	�4���P������R�����P�$�����P�R����������舿���������}����������r���3��3�_^[��`  ;��ޫ����]���������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   ������EP�M�蔵���EP�M�������E�P�M�|����M��p����ER��P���膖��XZ_^[���   ;��Ϊ����]Ë�   ������   ��s ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;��K�����E�P�MQ��*�B�H�у�;��)����E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M��_���P�M�艨���E�_^[���   ;�蝩����]� ���������������������������U����   SVWQ��4����3   ������Y�M���*�P��M��B<��;��@���_^[���   ;��0�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M��BL��;�迨��_^[���   ;�诨����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M��e����E�� L��E�_^[���   ;��E�����]����������������������U����   SVWQ��4����3   ������Y�M��M��0����E��t�E�P�ܓ�����E�_^[���   ;��ڧ����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� L��E���P�V������M������_^[���   ;��i�����]��������������������������U���T  SVWQ�������  ������Y�M��E�   j j h'  �M�脝���E�j h������������j ������Pj jjj �M�������������V���j jh�  j8h�  �M�蒘���M������j h��������走��j ������Pj jjj �M�袑��������� ���j j j j8h�  �M��1����M������M��ߡ���M��ס����l����̡���E�Ph'  �Ӵ�����E�Ph(  �´�����E�Ph2  豴������l���Ph�  蝴����j h��������� ���j h�����������h�  ��p����ʥ��������Ph'  ������Q������P�����Rh'  �\�����P��(���P蕶����P��@���Q腶����P��X���R�u�����Pj ��p���P�M��í����X����и����@����Ÿ����(���躸��������诸�������褸��������虸��j h������������j h������������h�  ���������������Ph�  ������Q������P������Rh'  �t�����P������P譵����P������Q蝵����P������R荵����Pj�����P�M��۬�������������������ݷ���������ҷ���������Ƿ��������輷��������豷��j h���� ����0���j h����P�������h�  ������������� ���Ph�����8���Q������P��P���Rh'  茊����P��h���P�Ŵ����P������Q赴����P������R襴����Pj������P�M������������ ����������������h���������8����߶����P����Զ���� ����ɶ��j h���������H���j h���������6���h�  ��P�������������P�M�Q������R�i�����P������Ph'  襉����P�����Q�޳����P�� ���R�γ����P��8���P辳����Pj��P���Q�M�������8��������� ������������������������������������������������M�蘶��j h����`����Y���j ��`���Pj jjj �M��F�����`���褵����P���腈��jhrdrb��P�������jhttub��P����/���j h|���x����������P���PjPjPj ��x���QhD h'  �M��*����U��B��x����,���j h ���E��H�|�����P���腊���M��ŵ���E�R��P�������XZ_^[��T  ;��e�����]Ð   �����   S�����   N�����   I�l���   D�P���   @�bbc dat4 dat3 dat2 dat1 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVW��(����6   �������EP��,���Q��*�B�H(�у�;�虞��P�M������,��������E_^[���   ;��r�����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P0��;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P4��;�臝��_^[���   ;��w�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E�_^[��]� �������������������������������U���$  SVWQ�������I   ������Y�M��M��\�����u3��  h'  ������衜��j j ������P�M�蜎��h'  �������~���j j �����$�����$haerf�����$������$������$�����$������P�M��č��h'  �� �������h���h  �j jh���h  �h'  �� ���P�M��|���j h������������h�  ��(����Л��j j �����P��(���Q�M�����������.����   _^[��$  ;�蛛����]��������������������������������������������������������������������������������������������U���  SVWQ��x�����   ������Y�M�葪���E�M�������M�胖���M��������7����E̍M��Ӂ�����Q����EЍE�Ph ���f������E��E��E��@   j havem�M蒗���E�j havem�M耗���E�j havem�M�n����E�j havem�M�\����E�j havem�M�J�����x���j havem�M�5�����l����E��x�����x���'  1��x���'  tJ��x����  ��  ��x���'  �Z  �  ��x���'  ��   ��x���'  ��   �\  j h���������ܣ��������P��������������1����E�P������Q�ס����P�Ԫ�����������
����E�P������Q谡����P譪���������������E�Ph ����������u,j h���������M���������P�l�����������袬���  j h������������������P�;������������q����k  �}�'  u,j h|�����������������P�������������7����}�'  u,j h`������譢�������P�̩���������������   �}� u,j h|���(����v�����(���P蕩������(����˫���}�u,j h`���@����D�����@���P�c�������@���虫����x���u,j hD���X���������X���P�.�������X����d�����l���u,j h(���p����ڡ����p���P���������p����/����,j h�������謡��������P�˨��������������j ������ǅ����   �M�谣��������R��P�$�����XZ_^[�Ĉ  ;��@�����]� ��   ,����   J����   Didata myicon �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;�贕��_^[���   ;�褕����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;��;���_^[���   ;��+�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;��˔��_^[���   ;�軔����]����������������������������U����  SVWQ��<����q   ������Y�M��M������M蔂����<�����<���NPIbt�F  j hvdpi�M�(���=byek�,  ��D���讚��Phcsak�E�P�M������D���莧���E�P�A�����j h����h���������h���P�M��w}����\�����h����P�����\��� ��   �M��>���h�  ������訓���E�P������Q�M��ը���M��8����E��E�    j h��������腝��j��E�P������Q�M������E��������Ѧ���E�+E�P�M���Q��t���R�M�������t���P�M��Ш����t���蚦���M�蒦���M�芦���E�P�=������EP�MQ�M������������M��`���������R��P��	�s~��XZ_^[���  ;�軒����]� �   �	����   �	����   �	����   �	����   �	t���   �	lw pos text input lastWord ���������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��*�B�H�у�;��w����E�_^[���   ;��d�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;�������E�_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M��EP�M��[x�������_^[���   ;�膐����]� ��������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bx��;��+���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M��BD��;�贏��_^[���   ;�褏����]� ����������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R��*�P�M��BP��;��1���P�M誙���� ���蛢���E_^[���   ;��
�����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M��B ��;�蠎��_^[���   ;�萎����]���������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R��*�P�M����   ��;�����P�M藘���� ���舡���E_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M��|��j h�   h,  j�j�hFB j�M����Or��_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M��EPj hFB �M���蒈��_^[���   ;�背����]� ���������������������������������U����  SVW������   ������h���������r��h����0����r�������P��0���Q��T���R�ա����P��x���P� �����P�M�Q��������x����2y����T����'y����0����y��������y���M�衋��j j��E�P�M��r������q����t%ǅ����    �M��˗���M���x���������  jj j j j �M��}��Ph ���K�����j hp��M��O���h��8��
Ph�/j�͓���������������� t�������5���������
ǅ���    j h�������������j h�����������������Q�U�R������P�������Px��������Pj ������QhFB ���������������������������������������������M������M�誖���M��w��������R��P�0��u��XZ_^[���  ;��2�����]Ë�   8����   e����   a����   \Help bmp fn ������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��M�耞���E�� ���M���芀���E�_^[���   ;�躈����]���������������������������U����   SVWQ��4����3   ������Y�M��M��z���E��t�E�P�Lt�����E�_^[���   ;��J�����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E�� ���E�_^[���   ;�������]����������������������U����   SVWQ��4����3   ������Y�M��M����͙���M��ϙ��_^[���   ;�膇����]�����������������������U����   SVWQ��4����3   ������Y�M��M��x��_^[���   ;��1�����]������������������U����   SVWQ��4����3   ������Y�M��M��*����E��t�E�P��r�����E�_^[���   ;��ʆ����]� ������������������������U����   SVWQ��4����3   ������Y�M��1p���M���E�_^[���   ;��l�����]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P��n�����E��     _^[���   ;�������]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M���j j���*�P�M��B��;��,����E�_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���j �EP��*�Q�M��B��;�蹄���E�_^[���   ;�覄����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EPj���*�Q�M��B��;��9����E�_^[���   ;��&�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��������]������������������U����   SVWQ��4����3   ������Y�M���*�P��M��B��;��p���_^[���   ;��`�����]���������������������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M�ow���E�_^[���   ;��������]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M����   ��;�葂��_^[���   ;�聂����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�H�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�H�у�;�藁�������_^[���   ;�老����]� ������������������������������U����   SVWQ��(����6   ������Y�M��EP�M������E�M��q��_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �BX�Ѓ�;�言��_^[���   ;�蘀����]�������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bt��;��;���_^[���   ;��+�����]� �������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M��
h��_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M��Bl��;��T��_^[���   ;��D����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M��g��_^[���   ;���~����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��[����E�EP�M�荑��_^[���   ;��^~����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*���   �H`�у�;���}��_^[���   ;���}����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;��x}��_^[���   ;��h}����]� ����������������������U����   SVWQ��(����6   ������Y�M���EP��*�Q�M����   ��;��}���E�}� u3���M�賀��_^[���   ;���|����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �B�Ѓ�;��x|��_^[���   ;��h|����]�������������������������U����   SVW��<����1   ������} t�E��<������*�b����<�����<���Q�UR�EP��r����_^[���   ;���{����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��k��_^[���   ;���z����]������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q��*�B<�H�у�;��cz���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����p��������
ǅ���    �E��@    _^[���   ;���y����]���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M���f���E��t�E�P�\e�����E�_^[���   ;��Zy����]� ������������������������U����   SVWQ������?   ������Y�M������P�ގ����P�M��rg�������������If�������_^[���   ;���x����]���������������������������U����   SVWQ��$����7   ������Y�M��E��x ufh ����Ph�/j��������,�����,��� t�MQ��,����E�����$����
ǅ$���    �U���$����B�E��x u3��Q�E��x t�E�3Ƀ8 �����9��EP��*�Q<��Ѓ�;���w���M���E��@   �E�3Ƀ8 ����_^[���   ;���w����]� �����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@   ��*�H<��Q��;��9w���M���E�3Ƀ8 ����_^[���   ;��w����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �4�E��x u3��'��E��HQ�U��P��*�Q<�B�Ѓ�;��v��_^[���   ;��uv����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u��*�H��#��EP�M��R��*�H<�Q�҃�;���u��_^[���   ;���u����]� ��������������������������������U����   SVW��@����0   �����󫹄*�Df��_^[���   ;��u����]���������������������U����   SVW��@����0   ������EP��*�3���_^[���   ;��0u����]�����������������U���  SVW�������B   ������EP��*����P�M��i��j h\ �������~��j �E�P�����Q�M��z�������������������&�����������t�M�{���M������E�9j�E�P�M���g��j�j��EP�M�Q�M��?s���E�P�M��~���M��Ї���ER��P�4(��_��XZ_^[��  ;��.t����]Ë�   <(����   X(����   T(str pos ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M��B@��;��ds��_^[���   ;��Ts����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��PH��;���r��_^[���   ;���r����]� �������������������������������������U���,  SVW�������K   ������EP��*�s���P�M���|��j h\ �������t|��j �E�P������Q�M��6x�������������������超����������t�M�x���M�蛅���E�   j�E�P�M��xe��j�j��EP�M�Q�M���p��j h\ �������{��j �E�P�����Q�M��w�������������������2�����������t�M�"x���M������E�9j�E�P�M���d��j�j��EP�M�Q�M��Kp���E�P�M��{���M��܄���ER��P�(+��\��XZ_^[��,  ;��:q����]Ë�   0+����   L+����   H+str pos ����������������������������������������������������������������������������������������������������������������U���P  SVW�������T   ������EP��*�c���P�M���z��j h\ �������dz��j �E�P������Q�M��&v�������������������覃����������t�M�v���M�苃���E�>  j�E�P�M��hc��j�j��EP�M�Q�M��n��j h\ ��������y��j �E�P������Q�M��u��������������������"�����������t�M�v���M������E�   j�E�P�M���b��j�j��EP�M�Q�M��8n��j h\ ������\y��j �E�P�����Q�M��u������������������螂����������t�M�u���M�胂���E�9j�E�P�M��cb��j�j��EP�M�Q�M��m���E�P�M�Ty���M��H����ER��P��-�^Z��XZ_^[��P  ;��n����]Ë�   �-����   �-����   �-str pos ��������������������������������������������������������������������������������������������������������������������������������������������U���t  SVW�������]   ������EP��*���P�M��9x��j h\ �������w��j �E�P������Q�M��vs��������������������������������t�M��s���M��ۀ���E��  j�E�P�M��`��j�j��EP�M�Q�M��l��j h\ �������0w��j �E�P������Q�M���r��������������������r�����������t�M�bs���M��W����E�>  j�E�P�M��4`��j�j��EP�M�Q�M��k��j h\ �������v��j �E�P������Q�M��nr�������������������������������t�M��r���M������E�   j�E�P�M��_��j�j��EP�M�Q�M��k��j h\ ������(v��j �E�P�����Q�M���q�������������������j����������t�M�Zr���M��O���E�9j�E�P�M��/_��j�j��EP�M�Q�M��j���E�P�M� v���M�����ER��P��0�*W��XZ_^[��t  ;��rk����]Ë�   �0����   1����   1str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������EP��*�Q<�B�Ѓ�;��Pj��_^[���   ;��@j����]���������������������������������U���p  SVW�������\   ������ǅ����    j h����������s��P�S�����E��������I}���}� u3���   �E�    �E�P�M���X���E�P�M�Q�M���i������   �}���   �M���W���E��}� tF�EP��������o��������Pj������Q�M��Rq������������R����tǅ����   �
ǅ����    ��������������������t��������������}|����������t��������������`|����������t�EԉE�������E�R��P��3�^T��XZ_^[��p  ;��h����]Ë�   �3����   �3����   �3����   �3browse dat id ��������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �BT�Ѓ�;��g��_^[���   ;��g����]�������������������������U���d  SVW�������Y   ������ǅ����    �} u6j h���������Kq��P�Q�����E�������z���} u3��$  �E�    �EP�M��HV���E�P�M�Q�M��Jg������   �}���   �M��GU���Eă}� tF�EP�������Dm��������Pj������Q�M��n�����������0P����tǅ����   �
ǅ����    ��������������������t���������������y����������t��������������y����������t�E��E��2�+�}�u%�}� t�EP�M���y�����O����t�E��E��������E�R��P��6�Q��XZ_^[��d  ;���e����]ÍI    �6����   �6����   �6����   �6browse dat id ��������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �BH�Ѓ�;���d��_^[���   ;��d����]�������������������������U����   SVW������:   ������} u3��   �EP�M��S���E�    �E�    �E�P�M�Q�M��d����tT�}�t�}�u"�EP�M��R��P�T������t�   �*�$�}�u�EP�M���w�����M����t�   ��3�R��P��8�O��XZ_^[���   ;���c����]�   �8����   �8����   �8����   �8dat id browse ����������������������������������������������������������������������������������U����   SVW��@����0   �����󫡘*�H<��Q��;��c��_^[���   ;���b����]�������������������������U����   SVW��@����0   ������E��*��*� _^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M���h����E�P��*�Q$�BD�Ѓ�;��Cb���E�_^[���   ;��0b����]���������������������������������U����   SVWQ��4����3   ������Y�M��M��bh����E�P��*�Q$�BD�Ѓ�;���a����EP�M�Q��*�B$�Hd�у�;��a���E�_^[���   ;��a����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��g����E�P��*�Q$�BD�Ѓ�;��a����EP�M�Q��*�B$�H�у�;���`���E�_^[���   ;���`����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��g����E�P��*�Q$�BD�Ѓ�;��c`����E�P�MQ��*�B$�HL�у�;��A`���E�_^[���   ;��.`����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q$�BH�Ѓ�;��_���M��1s��_^[���   ;��_����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�HL�у�;��7_��_^[���   ;��'_����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q$�M��B��;��^��_^[���   ;��^����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q$�M��Bl��;��;^��_^[���   ;��+^����]� �������������������������U����   SVWQ��4����3   ������Y�M���*�P$��M��Bp��;���]��_^[���   ;���]����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q$�B�Ѓ�;��[]��_^[���   ;��K]����]����������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q��*�B$�H�у�;���\��P�M�]g���� ����Np���E_^[���   ;��\����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H�у�;��G\��_^[���   ;��7\����]� �������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q��*�B$�H �у�;���[��P�M�f��������	I���E_^[���   ;��[����]� �������������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q��*�B$�H$�у�;��$[��P�M�f��������iH���E_^[���   ;���Z����]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M��eO�����B���������G���E_^[���   ;��qZ����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q$�B(�Ѓ�;��Z��_^[���   ;���Y����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q$�Bh�Ѓ�;��Y��_^[���   ;��Y����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H,�у�;��'Y��_^[���   ;��Y����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H0�у�;��X��_^[���   ;��X����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H4�у�;��'X��_^[���   ;��X����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H8�у�;��W��_^[���   ;��W����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��*�B$�HL�у�;��'W���E�_^[���   ;��W����]� ����������������������������������U����   SVW������9   ������EP�M��a����EP�M�Q��*�B$�H@�у�;��V���E�P�M�a���M���C���ER��P��E� B��XZ_^[���   ;��hV����]�    F����   Ffn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H@�у�;���U���E�_^[���   ;���U����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H<�у�;��WU��_^[���   ;��GU����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�H<�у�;���T�������_^[���   ;���T����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H$�QP�҃�;��TT��_^[���   ;��DT����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B$�HT�у�;���S��_^[���   ;���S����]� �������������������������������������U����   SVW��@����0   �����󫡘*�H$��QX��;��hS��_^[���   ;��XS����]�������������������������U����   SVW��@����0   �������EP��*�Q$�B\�Ѓ�;�� S��_^[���   ;���R����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q$�B`�Ѓ�;��R��_^[���   ;��oR����]� �����������������������������U����   SVW��@����0   �����󫡘*�H(����;��R��_^[���   ;��	R����]��������������������������U����   SVW��@����0   �������E�Q��*�B(�H�у�;��Q���E�     _^[���   ;��Q����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR��*�P(�M��B��;��Q��_^[���   ;��Q����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���*�P(��M��B��;��P��_^[���   ;��P����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��B��;��+P��_^[���   ;��P����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P(�M��B��;��O��_^[���   ;��O����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B(�M��P ��;��7O��_^[���   ;��'O����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ��*�B(�M��P��;��N��_^[���   ;��N����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P(�M��B$��;��4N��_^[���   ;��$N����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���*�P(��M��B(��;���M��_^[���   ;��M����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P(��M��B,��;��PM��_^[���   ;��@M����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P(��M��B0��;���L��_^[���   ;���L����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��B4��;��kL��_^[���   ;��[L����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��BX��;���K��_^[���   ;���K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��B\��;��K��_^[���   ;��{K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��B`��;��K��_^[���   ;��K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bd��;��J��_^[���   ;��J����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bh��;��;J��_^[���   ;��+J����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bx��;���I��_^[���   ;��I����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bl��;��[I��_^[���   ;��KI����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bt��;���H��_^[���   ;���H����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��Bp��;��{H��_^[���   ;��kH����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M���9����t2�M��Q�M���9����t�U��R�M��9����tǅ0���   �
ǅ0���    ��0���_^[���   ;���G����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��S����t8�MQ�A�$�M��S����t"�UQ�B�$�M��{S����tǅ0���   �
ǅ0���    ��0���_^[���   ;��G����]� ������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M���E����t2�M��Q�M���E����t�U��R�M���E����tǅ0���   �
ǅ0���    ��0���_^[���   ;��WF����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M���4����t<�M���A�$�M���4����t$�U���B�$�M��4����tǅ0���   �
ǅ0���    ��0���_^[���   ;��E����]� ����������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��B?����tE�M��Q�M��/?����t2�U��R�M��?����t�E��$P�M��	?����tǅ0���   �
ǅ0���    ��0���_^[���   ;���D����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��Q<����tE�M��Q�M��><����t2�U��R�M��+<����t�E��$P�M��<����tǅ0���   �
ǅ0���    ��0���_^[���   ;���C����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M���(����tE�M��Q�M���(����t2�U��0R�M���(����t�E��HP�M��(����tǅ0���   �
ǅ0���    ��0���_^[���   ;��$C����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M���O����tE�M��Q�M��O����t2�U��0R�M��O����t�E��HP�M��O����tǅ0���   �
ǅ0���    ��0���_^[���   ;��TB����]� ��������������������������������������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M��X(����u3���   �}� u)������DH��P�M�cW��������-U���   �   ��h` ����P�M�Q��*�B���   �у�;��vA���E��}� uj��M��B��3��Lj �E�P�M�Q�M��T����u�E�P�8����3��&j �E��P�M�Q�M�TC���E�P��7�����   R��P�p[�,��XZ_^[���   ;���@����]�    x[����   �[����   �[c len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q�B�Ѓ�;��@��_^[���   ;��@����]� �����������������������������U����   SVWQ������?   ������Y�M��M��BF���E�P�M��Y7����uǅ���    �M��S��������$�E�P�M�D'��ǅ���   �M���R�������R��P�]�
+��XZ_^[���   ;��R?����]�    ]����   $]str ��������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�P�M���.����u3���E�����؋M��   R��P��]�H*��XZ_^[���   ;��>����]� ��   �]����   �]c ��������������������������������������U����   SVWQ��4����3   ������Y�M��} ����Q�M��ZJ��_^[���   ;��>����]� ��������������������U����   SVWQ������=   ������Y�M�j �M��3�����E���h` ����P�M�Q��*�B���   �у�;��=���Eԃ}� uj��M��>��3��dj �E�P�M�Q�M�B���E�P�M��,R����t �M�Q�U�R�M��8F����tǅ���   �
ǅ���    ������E�E�P��3�����E�R��P�t_�(��XZ_^[���   ;���<����]�    |_����   �_mem ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bd��;��;<��_^[���   ;��+<����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P�M��Bh��;���;��_^[���   ;��;����]� ����������������������������������U����   SVWQ������<   ������Y�M��� ���P�M�Y#��P�M��I��������� ����N�������_^[���   ;��*;����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q(�M��B8��;��:��_^[���   ;��:����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q(�M��B<��;��J:��_^[���   ;��::����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q(�M��B@��;���9��_^[���   ;���9����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q(�M��BD��;��j9��_^[���   ;��Z9����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��BH��;���8��_^[���   ;���8����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B(�M��P|��;��8��_^[���   ;��w8����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q(�M��BL��;��8��_^[���   ;���7����]� �������������������������U����   SVWQ��4����3   ������Y�M�����E�$��*�P(�M��BT��;��7��_^[���   ;��7����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$��*�P(�M��BP��;��7��_^[���   ;��	7����]� �����������������������U����   SVW��@����0   �����󫡘*�H(��Q��;��6��_^[���   ;��6����]�������������������������U����   SVW��@����0   �������E�Q��*�B(�H�у�;��N6���E�     _^[���   ;��56����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP��*�Q(�M����   ��;��5��_^[���   ;��5����]�( ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��*�B(�H�у�;�� 5��_^[���   ;��5����]���������������������������������U����   SVW��@����0   �����󫡘*�H,��Q,��;��4��_^[���   ;��4����]�������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B4��;��P4��_^[���   ;��@4����]���������������������������������U����   SVW��@����0   �������E�Q��*�B,�H0�у�;���3���E�     _^[���   ;���3����]��������������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B8��;��`3��_^[���   ;��P3����]���������������������������������U����   SVWQ������<   ������Y�M������P��*�Q,�M��B<��;���2��P�M��=��������- ���E_^[���   ;���2����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q��*�B,�M��P@��;��T2��P�M��<���� ����E���E_^[���   ;��-2����]� �������������������������������������������U����   SVW��@����0   �������j j ��*�H,��҃�;���1��_^[���   ;��1����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H,�Q�҃�;��D1��_^[���   ;��41����]� ����������������������������������U����   SVW��@����0   �������E�Q��*�B,�H�у�;���0���E�     _^[���   ;��0����]��������������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B��;��P0��_^[���   ;��@0����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B��;���/��_^[���   ;���/����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B��;��p/��_^[���   ;��`/����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B ��;�� /��_^[���   ;���.����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B$��;��.��_^[���   ;��.����]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P,��M��B(��;�� .��_^[���   ;��.����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B,�M��P��;��-��_^[���   ;��-����]� �������������������������������������U����   SVWQ������<   ������Y�M������P��*�Q,�M��B��;��(-��P�M�8��������m���E_^[���   ;��-����]� �������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��D  �҃�;��,��_^[���   ;��,����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��H  �҃�;��&,��_^[���   ;��,����]�����������������������U����   SVW��@����0   �������EP��*�Q��L  �Ѓ�;��+��_^[���   ;��+����]������������������������������U����   SVW��@����0   �������EP�MQ��*�B�H�у�;��L+��_^[���   ;��<+����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H�Q�҃�;���*��_^[���   ;���*����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B�H�у�;��l*��_^[���   ;��\*����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H�Q�҃�;���)��_^[���   ;���)����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B�H�у�;��)��_^[���   ;��|)����]�����������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;��)��_^[���   ;��	)����]��������������������������U����   SVW��@����0   �������EP��*�Q�B�Ѓ�;��(��_^[���   ;��(����]���������������������������������U���  SVW�������E   ������E�P�M�R���M�������uǅ����    �M�����������   j�E�P�S������u*�E�P�:.������uǅ����    �M��N���������Tj�EP�������u*�EP�,������uǅ���    �M����������ǅ���   �M����������R��P��t�0��XZ_^[��  ;��x'����]�   �t����   �tparent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP��*�Q�B �Ѓ�;���&��_^[���   ;���&����]���������������������������������U����   SVW��@����0   �������EP�MQ��*�B�H(�у�;��\&��_^[���   ;��L&����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��*�B��  �у�;���%��_^[���   ;���%����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q��   �Ѓ�;��a%��_^[���   ;��Q%����]����������������������������������U����   SVW��@����0   �������EP��*�Q��  �Ѓ�;���$��_^[���   ;���$����]������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��  �҃�;��v$��_^[���   ;��f$����]�����������������������U����   SVW������9   ������� ���P��*�Q�B$�Ѓ�;��$��P�M��.���� ����R���E_^[���   ;���#����]���������������������������������������U����   SVW������9   ������� ���P��*�Q���  �Ѓ�;��z#��P�M�a.���� �������E_^[���   ;��S#����]������������������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;���"��_^[���   ;���"����]��������������������������U���$  SVW�������I   ������ǅ8���    �=p/ t!������P�p/�y����8�����������������*����8���������������������������R�M�'-����8�����t��8����������s����8�����t��8�����������V���E_^[��$  ;���!����]�����������������������������������������������������������U����   SVW������9   �������EP�� ���Q��*�B���  �у�;��f!��P�M�M,���� �������E_^[���   ;��?!����]��������������������������������U����   SVW��@����0   ������j�EP�p&�����E_^[���   ;��� ����]������������������������������U����   SVW��@����0   �����󫡘*�H���   ��;�� ��_^[���   ;��u ����]����������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;�� ���E�     _^[���   ;�� ����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M����;����_^[���   ;������]� ������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M��B��;�� ��_^[���   ;������]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B`��;��;��_^[���   ;��+����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bd��;�����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bh��;��[��_^[���   ;��K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bl��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bp��;��{��_^[���   ;��k����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bt��;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��Bx��;��+��_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B|��;��K��_^[���   ;��;����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;��h��_^[���   ;��X����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;��x����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;��8��_^[���   ;��(����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;��X��_^[���   ;��H����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B��  �у�;��t��_^[���   ;��d����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��t��_^[���   ;��d����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q��*�B �H$�у�;������tǅ0���   �
ǅ0���    ��0���_^[���   ;��Q����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR��*�H �QL�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q��*�B �H(�у�;��M���   _^[���   ;��8����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q�M��B��;�����_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q�M��B��;��Z��_^[���   ;��J����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q�M��B��;�����_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP��*�Q�M��B��;��z��_^[���   ;��j����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B��;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P\��;��'��_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$��*�P�M��B ��;����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$��*�P�M��B$��;��)��_^[���   ;������]� �����������������������U����   SVWQ��4����3   ������Y�M�����E�$��*�P�M��B(��;����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B,��;��;��_^[���   ;��+����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B0��;�����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B4��;��[��_^[���   ;��K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B8��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B<��;��{��_^[���   ;��k����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B@��;����_^[���   ;���
����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BD��;��
��_^[���   ;��
����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BH��;��+
��_^[���   ;��
����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BL��;��	��_^[���   ;��	����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BP��;��K	��_^[���   ;��;	����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M����   ��;�����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BT��;��[��_^[���   ;��K����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B��  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M����   ��;��\��_^[���   ;��L����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M����   ��;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��PX��;��g��_^[���   ;��W����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;��x��_^[���   ;��h����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��$��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��4��_^[���   ;��$����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;��M��_^[���   ;��=����]������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M����   ��;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��*�B���   �у�;��]��_^[���   ;��M����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q��   �Ѓ�;��� ��_^[���   ;��� ����]����������������������������������U����   SVW��(����6   �������EP�MQ��,���R��*�H���  �҃�;��c ��P�M��
����,��������E_^[���   ;��< ����]���������������������������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;������_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B8�HD�у�;��W���_^[���   ;��G�����]� �������������������������������������U����   SVW��@����0   �����󫡘*�H8��Q<��;������_^[���   ;��������]�������������������������U����   SVW��@����0   �������E�Q��*�B8�H@�у�;��~����E�     _^[���   ;��e�����]��������������������������������������U����   SVW��@����0   �����󫡘*�H8����;��	���_^[���   ;��������]��������������������������U����   SVW��@����0   �������E�Q��*�B8�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q8�B�Ѓ�;�����_^[���   ;��������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H8�Q�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q8�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B8�H �у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�H8�Q$�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P��*�Q8�B�Ѓ�;�����_^[���   ;��s�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H8�Q(�҃�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q8�B,�Ѓ�;�����_^[���   ;��o�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q8�B�Ѓ�;������_^[���   ;��������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�H8�Q�҃�;��x���_^[���   ;��h�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H8�Q0�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q8�B4�Ѓ�;��o���_^[���   ;��_�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B8�H8�у�;������_^[���   ;��������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q��x  �Ѓ�;��q���_^[���   ;��a�����]����������������������������������U����   SVW��@����0   �������EP�MQ��*�B��|  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;�����_^[���   ;��y�����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;�����_^[���   ;��	�����]��������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��*�Q�B,�Ѓ�;��@���_^[���   ;��0�����]���������������������������������U����   SVW��(����6   ������M��g�����E�P��*�Q�B8�Ѓ�;�������E�P�M�>����M��2���ER��P�Ш�H���XZ_^[���   ;�������]�   ب����   �str ����������������������������������������U����   SVW��@����0   �����󫡘*�H��Q<��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ��*�B�H@�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �����󫡘*�H��QD��;��H���_^[���   ;��8�����]�������������������������U����   SVW��@����0   �����󫡘*�H��QH��;������_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H�QL�҃�;��y���_^[���   ;��i�����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B�HP�у�;�����_^[���   ;��������]�����������������������������U����   SVW��@����0   �������EP��*�Q��<  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��*�Q��,  �Ѓ�;��-���_^[���   ;�������]������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP��*�Q���   �Ѓ�;�����_^[���   ;�������]���������������������������������������U����   SVW��@����0   �����󫡘*�H�􋑼   ��;��%���_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡘*�H���  ��;������_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�.  ��*�B���   �у�;��H���_^[���   ;��8�����]�����������������������������������������U����   SVW��@����0   �������EP��*�Q�B�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP��*�Q��\  �Ѓ�;��]���_^[���   ;��M�����]������������������������������U����   SVW������<   ������EPj h� ���������P�M�Q�������������^ ����E�P��*�Q�B�Ѓ�;�������M��8 ��R��P�ȯ�Q���XZ_^[���   ;�������]Ð   Я����   ܯs ��������������������������������������������������U����   SVW��@����0   �������EP��*�Q�BT�Ѓ�;�����_^[���   ;�� �����]���������������������������������U����   SVW��@����0   �������EP��*�Q�BX�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP��*�Q�B\�Ѓ�;��0���_^[���   ;�� �����]���������������������������������U����   SVW��@����0   �����󫡘*�H��Q`��;������_^[���   ;�������]�������������������������U����   SVW��@����0   �����󫡘*�H��Qd��;��h���_^[���   ;��X�����]�������������������������U����   SVW��@����0   �����󫡘*�H��Qh��;�����_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP��*�Q�Bl�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP��*�Q�Bp�Ѓ�;��0���_^[���   ;�� �����]���������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H�Qt�҃�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��*�Q��D  �Ѓ�;��M���_^[���   ;��=�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q��  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ��*�B�Hx�у�;��\���_^[���   ;��L�����]�����������������������������U����   SVW��@����0   �������EP�MQ��*�B��@  �у�;������_^[���   ;��������]��������������������������U����   SVW������9   ������M�������E�P�MQ��*�B�H|�у�;��t����E�P�M�X����M������ER��P�$������XZ_^[���   ;��<�����]�   ,�����   8�fn �����������������������������������������������������U����   SVW��@����0   �������EP�MQ��*�B���   �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ��*�B��h  �у�;��9���_^[���   ;��)�����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q��d  �Ѓ�;������_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;��F���_^[���   ;��6�����]�����������������������U����   SVW��@����0   �����󫡘*�H�􋑄   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ��*�B��l  �у�;��y���_^[���   ;��i�����]��������������������������U����   SVW��@����0   �������EP��*�Q��   �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��$����7   ������M�������E�P��*�Q���   �Ѓ�;��%����E�P�M�����M������ER��P�t�����XZ_^[���   ;��������]Ð   |�����   ��bc �����������������������������������������������������U����   SVW��@����0   �����󫡘*�H��`  ��;��e���_^[���   ;��U�����]����������������������U����   SVW��@����0   �������EP��*�Q��  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW�� ����8   �������EP��$���Q��*�B���   �у�;������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��N�����]�����������������������������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ��*�B���   �у�;��W���_^[���   ;��G�����]����������������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���   �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���   �҃�;��f���_^[���   ;��V�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;�����_^[���   ;��v�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���   �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ��*�B���   �у�;��9���_^[���   ;��)�����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B���   �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;��]���_^[���   ;��M�����]������������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;��}���_^[���   ;��m�����]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��*�Q���   �Ѓ�;��������u3���E�R��P�������XZ_^[���   ;��������]�   ������   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��*�Q���   �Ѓ�;�������u3���E�R��P�������XZ_^[���   ;��������]�   ������   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P��*�Q���   �Ѓ�;�������u3���E�R��P�p�����XZ_^[���   ;��������]�   x�����   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP��*�Q��8  �Ѓ�;��=���_^[���   ;��-�����]������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�����P�U�R��*�H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�J���P�U�R��*�H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P��*�Q0���   �Ѓ�(;������_^[���   ;�������]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B0���   �у�;��8���_^[���   ;��(�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q0���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H0���   �҃�;��A���_^[���   ;��1�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B0���   �у�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q0���   �Ѓ�;��8���_^[���   ;��(�����]�������������������������U����   SVW��@����0   �����󫡘*�H0�􋑤   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������E�Q��*�B0���   �у�;��k����E�     _^[���   ;��R�����]�����������������������������������U����   SVW��@����0   �������EP��*�Q��H  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��*�Q��T  �Ѓ�;��}���_^[���   ;��m�����]������������������������������U����   SVW��@����0   �����󫡘*�H��p  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡘*�H���  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��M���_^[���   ;��=�����]������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��m���_^[���   ;��]�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q���  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��*�B���  �у�;��m���_^[���   ;��]�����]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P��*�Q��X  �Ѓ�;������P�M�5�����,��������E_^[���   ;��������]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q��*���   �H�у�;��?����E�_^[���   ;��,�����]� ������������������������������������������U����   SVW������=   ������j hLGOg�����蜺��PhicMC�E�P�����������裴���M�������u�M�����M��Q����E��M�����P�M�����M��3����ER��P���	���XZ_^[���   ;��Q�����]Ð   �����   $�dat ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ��*�B��  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP��*�Q��\  �Ѓ�;��M���_^[���   ;��=�����]������������������������������U����   SVW������9   ������EP��MQ�� ���R��*�H��t  �҃�;���������˱���� ��������E_^[���   ;�������]�������������������������������U����   SVW��(����6   �������EP��,���Q��*�B���  �у�;��F���P�M������,��������E_^[���   ;�������]��������������������������������U����   SVW��(����6   �������EP��,���Q��*�B���  �у�;�����P�M�/�����,���� ����E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��-���_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��M���_^[���   ;��=�����]������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ��*�B���  �у� ;������_^[���   ;�������]����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR��*�H���  �҃�$;��.���_^[���   ;�������]�������������������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q��*�B��t  �у�;�����P�M�!�����,��������E_^[���   ;�������]����������������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q��*�B���  �у�;��
���P�M�Q�����,��������E_^[���   ;��������]������������������������������������U����   SVW��@����0   �������EP��*�Q��8  �Ѓ�;��}���_^[���   ;��m�����]������������������������������U����  SVW��(����6  ������h3ŉE��E�E�E�P�MQh   ������R�������������Ph� ��*�Q��4  �Ѓ�;�������E�    R��P����i���XZ_^[�M�3��������  ;�������]ÍI    ������   ��t ��������������������������������������������������������������U����   SVW��4����3   ������} 3��^�EP�MQ�UR�EP茾�����E��}� |�E��9E�|/�}� }h� ����P蒫�����EE�@� �E���E��E�_^[���   ;�������]���������������������������������������U����   SVW��@����0   �������EP�MQ��*�B��0  �у�;��I���_^[���   ;��9�����]��������������������������U����   SVW��(����6   �������,���P��*�Q��  �Ѓ�;������P�M�S�����,����D����E_^[���   ;�������]������������������������������������U����   SVW��(����6   �������,���P��*�Q��  �Ѓ�;��J���P�M�������,��������E_^[���   ;��#�����]������������������������������������U����   SVW������=   �������T�����u�\h���M�薯���EPh���M�躻���EPh���M�詻��j �E�PhicMC�����Q�y�����������=����M��k���R��P������XZ_^[���   ;��V�����]Ë�   �����    �msg ������������������������������������������������������������U����   SVW������=   �������T�����u�M�N����E�^h!���M�苮���EPh!���M�诺��j �E�PhicMC�����Q���������p���P�M����������3����M��a����ER��P������XZ_^[���   ;��I�����]Ð    �����   ,�msg ����������������������������������������������������������������U����   SVW������=   �������D�����u�M�>����E�^h����M��{����EPh����M�蟹��j �E�PhicMC�����Q�o��������`���P�M�����������#����M��Q����ER��P�(�����XZ_^[���   ;��9�����]Ð   0�����   <�msg ����������������������������������������������������������������U���   SVW�� ����@   �������4�����u3��^h#���M��t����EPh#���M�蘸��j �E�PhicMC�����Q�h���������������������������M��M��������R��P�0�����XZ_^[��   ;��2�����]Ë�   8�����   D�msg ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �B8�Ѓ�;�蘼��_^[���   ;�舼����]�������������������������U���   SVW�� ����@   �������������u3��^hs���M������EPhs���M��(���j �E�PhicMC�����Q����������\������������������M��ݤ�������R��P����z���XZ_^[��   ;��»����]Ë�   ������   ��msg ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��*�H���  �҃�;�����_^[���   ;��
�����]���������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��@  �҃�;�覺��_^[���   ;�薺����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��*�H���  �҃�;��*���_^[���   ;�������]���������������������������U����   SVW��@����0   ������E�8 t#��E�Q��*�B��D  �у�;�賹���E�     _^[���   ;�蚹����]���������������������������U����   SVW��@����0   �������EP��*�Q��H  �Ѓ�;��=���_^[���   ;��-�����]������������������������������U����   SVW��@����0   �������EP��*�Q��L  �Ѓ�;��͸��_^[���   ;�轸����]������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��P  �҃�;��V���_^[���   ;��F�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��T  �҃�;�����_^[���   ;��ַ����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��X  �҃�;��v���_^[���   ;��f�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H��\  �҃�;�����_^[���   ;��������]�����������������������U����   SVW��@����0   �����󫡘*�H��d  ��;�襶��_^[���   ;�蕶����]����������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP��*�Q��h  �Ѓ�;��%���_^[���   ;�������]��������������������������������������U����   SVW��@����0   �������EP�MQ��*�B��l  �у�;�詵��_^[���   ;�虵����]��������������������������U����   SVW��@����0   �����󫡘*�H�􋑄  ��;��E���_^[���   ;��5�����]����������������������U����   SVW��$����7   �������EP��(���Q��*�B���  �у�;��ִ��P�M�R�����(���趝���E_^[���   ;�说����]��������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��M���_^[���   ;��=�����]������������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��ݳ��_^[���   ;��ͳ����]������������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;��i���_^[���   ;��Y�����]��������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;�膲��_^[���   ;��v�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;�覱��_^[���   ;�薱����]�����������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;��=���_^[���   ;��-�����]������������������������������U����   SVW��@����0   �������EP�MQ��*�B��$  �у�;��ɰ��_^[���   ;�蹰����]��������������������������U����   SVW��@����0   �������EP��*�Q��(  �Ѓ�;��]���_^[���   ;��M�����]������������������������������U����   SVW��@����0   �������EP��*�Q��,  �Ѓ�;�����_^[���   ;��ݯ����]������������������������������U����   SVW��@����0   �����󫡘*�H��0  ��;�腯��_^[���   ;��u�����]����������������������U����   SVW��@����0   �����󫡘*�H��<  ��;��%���_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q���  �Ѓ�;�豮��_^[���   ;�衮����]����������������������������������U����   SVW��@����0   �����󫡘*�H���  ��;��E���_^[���   ;��5�����]����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;��֭��_^[���   ;��ƭ����]�����������������������U����   SVW��4����3   ������j �M�"����E��}� t�E�P譮�����E�P�8�����R��P� ������XZ_^[���   ;��B�����]Ë�   (�����   4�c ������������������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ��*�B��  �у� ;�衬��_^[���   ;�葬����]����������������������������������U����   SVW��@����0   �����󫡘*�H��P  ��;��5���_^[���   ;��%�����]����������������������U����   SVWQ��4����3   ������Y�M��E���P������_^[���   ;��ʫ����]���������������������������U����   SVW��@����0   �������EP��*���   ���   �Ѓ�;��j���_^[���   ;��Z�����]���������������������������U����   SVWQ������:   ������Y�M��M�<�������������NIVbb�����NIVb�  �����TCAb5�����TCAb��  �����$'  ��  �����MicM�.  ��  �����INIbt]�  �����atni-�����atnit6�����ckhc�Z  �����ytsdt\�  �����cnys��   �o  谙���e  �E��x t
�   �T  �E��@   �E����M��B��;������/  �E����M��B��;�������E��@    �  �E��x u
�   ��   �E����M��B��;�迩����   j hIicM�M萦���E��EP�M�Q�U���M��P��;�芩���   j hIicM�M�[����E��EP�M�Q�U���M��P��;��U����uj hdiem�M�)����E��EP�M�Q�U���M��P��;��#����E��E��=�E����M��B��;������%�!��EP�M���M��B��;������   �3�_^[���   ;��Ψ����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� ��E�Ph����*�Q0��Ѓ�;��Χ���M��A�E��@    �E�_^[���   ;�諧����]��������������������������������������������U���$  SVW�������I   �������E�    �M�蹍���} tg��EP��*�Q4�B�Ѓ�;��+����EЃ}� uǅ����    �M�������������   ��E�P�MQ�UЋ�MЋP(��;������E��b��EP��*�Q0�B�Ѓ�;��Ħ���Eă}� uǅ����    �M�蝏���������g��E�P�MQ�Uċ�MċP ��;�胦���E��M�裔�����t"��E�P�MQ��*�B0�Hx�у�;��Q����E��������M��4���������R��P�H��ё��XZ_^[��$  ;�������]Ð   P�����   \�result �������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�<������E�_^[���   ;��:�����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �E��x t!��E��HQ��*�B0�H�у�;��Ƥ���E��@    _^[���   ;�謤����]���������������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B0���   �у�;��5���_^[���   ;��%�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H0���   �҃�;�貣��_^[���   ;�袣����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��M��e�����P��*�H0���   �҃�;��4���_^[���   ;��$�����]�������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j4�E��HQ��*�B0���   �у�(;�裢��_^[���   ;�蓢����]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j;�E��HQ��*�B0���   �у�(;�����_^[���   ;�������]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�远��P��*�Q0���   �Ѓ�;�菡��_^[���   ;�������]� �����������������������������U���   SVWQ�� ����@   ������Y�M��E P�M�貞���EPh8kds�M��!����E�    ��E�P�M�Qj �UR�EP�MQ�UR�EPj2�M������P��*�Q0���   �Ѓ�(;��Ϡ���EЉ�����M�貉�������R��P����O���XZ_^[��   ;�藠����]� �   ������   ������   ��r customdata �����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������P��*�H0���   �҃�;��ԟ��_^[���   ;��ğ����]�������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��t��j j j j j �E Pj �MQj�U��BP��*�Q0���   �Ѓ�(;��2�����EP�MQ�UR�EPj �MQ�U��BP��*�Q0���   �Ѓ�;������_^[���   ;�������]� ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ��*�B0�H�у�;��[���_^[���   ;��K�����]����������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;�������]� �������������������������������U����   SVWQ������9   ������Y�M��E��x uj �M�����E�X�M������P�EP�M�Q���P�M��QR�� ���P��*�Q0���   �Ѓ�;��P���P�M藝���� ���������E_^[���   ;��)�����]� �������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H0�Q�҃�;��%���_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��x u�7��j j j j j j �EPj j�M��QR��*�H0���   �҃�(;�臛��_^[���   ;��w�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�p�����P�EP�M�ܑ��P�M��QR��*�H0�Q�҃�;�����_^[���   ;��֚����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�И����P�M�@���P�E��HQ��*�B0���   �у�;��F���_^[���   ;��6�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M�0�����P�EP�M蜐��P�M��QR��*�H0�Q\�҃�;�覙��_^[���   ;�薙����]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��_�E��ًU�
�E��ًU�
��EP�MQ�U��BP��*�Q4�Bh�Ѓ�;�������E�E��ًU�
�E��ًU�
�E�_^[���   ;��͘����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��*�Q4�Bh�Ѓ�;��C���_^[���   ;��3�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��*�Q4�Bp�Ѓ�;�賗��_^[���   ;�裗����]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��_�E��ًU�
�E��ًU�
��EP�MQ�U��BP��*�Q4�Bp�Ѓ�;������E�E��ًU�
�E��ًU�
�E�_^[���   ;��ݖ����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M�h���h  ��EPj 3Ƀ} ����Qj �UR�EP�M��ߝ��_^[���   ;��J�����]� ����������������������������������������U���  SVWQ�������C   ������Y�M�htniv�M�輄���EPhulav�M������hgnlfhtmrf�M��ΐ���EPhinim�M�轐���EPhixam�M�謐���EPhpets�M�蛐���EPhsirt�M�芐���}   �u	�}$���t"�E Ph2nim�M��g����E$Ph2xam�M��V����E�P�MQ�����R�M�賀����荤�������������������M��~��������R��P�p諀��XZ_^[��  ;�������]�  �   x����   �msg ����������������������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M�htlfv�M��������E�$hulav�M��Y{���E,Phtmrf�M��*������E�$hinim�M��2{�����E�$hixam�M��{�����E$�$hpets�M��{���EDPhsirt�M��׎���E0��������Dz�E8��������D{,���E0�$h2nim�M���z�����E8�$h2xam�M��z���E@Phdauq�M��~����E�P�MQ�����R�M���~����赢������������������M��6|��������R��P�H	��~��XZ_^[��  ;�������]�@ �   P	����   \	msg ������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP��*�Q�M��B,��;��R���_^[���   ;��B�����]� ��������������������������������U���<  SVWQ�������O   ������Y�M�hgnrs�M�輀���EP������袋��������Qj�M��ѥ�������������EP�������w���������Qj�M�覥���������T����E�P�MQ�����R�M���|�����Ҡ��������������%����M��Sz��������R��P�,��|��XZ_^[��<  ;��8�����]� ��   4����   @msg ����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��$���_^[���   ;�������]� ����������������������������������U���  SVWQ�������C   ������Y�M�hCITb�M��~���EPhCITb�M�趢���EPhsirt�M�蟊���EPhulav�M�莊���E�P�MQ�����R�M���z�����Ş������������������M��Fx��������R��P�8��z��XZ_^[��  ;��+�����]� �   @����   Lmsg ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P8��;�臎��_^[���   ;��w�����]� �������������������������������������U����   SVWQ������<   ������Y�M�j �EP�� ���Q�M�v��P�UR�M��9���������� ����t��������_^[���   ;��������]� ������������������������������U����   SVWQ��4����3   ������Y�M��E,Pj �����$�����$htemf���E$�$���E�$���E�$���E�$�MQ�M���~��_^[���   ;��>�����]�( ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E,Pj �����$�����$hrgdf���E$�$�.����$���E�$�����$���E�$�����$���E�$�MQ�M��~��_^[���   ;��v�����]�( ����������������������������������������������������U����   SVW��@����0   �������E�H�58_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E,Pj �����$�����$htcpf�E$�5X���$�E�5X���$�E�5X���$���E�$�MQ�M���|��_^[���   ;��\�����]�( ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��M�M�P�����P�E P���E�$���E�$�MQ�M要��P�U��BP��*�Q0�B(�Ѓ�$;�诊��_^[���   ;�蟊����]� ���������������������������������������������U����   SVWQ������9   ������Y�M��E��x u3��J�M萈����P�E�P�M�����P�M��QR��*�H0�Q,�҃�;������E�3��}� ���M��E�R��P���u��XZ_^[���   ;��щ����]� �I    �����   �val ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M蠇����P�EP�M����P�M��QR��*�H0�Q,�҃�;�����_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��6�M� �����P�EP�M�l��P�M��QR��*�H0�Q0�҃�;��v���_^[���   ;��f�����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M�������u3��;�E��P�MQ�M��d�����u3�� �E��P�MQ�M��I�����u3���   _^[���   ;�趇����]� ������������������������������������U���   SVWQ�� ����@   ������Y�M��E��x u3��   �E�    �M覅����P�E�P�M�~��P�M��QR��*�H0�Q8�҃�;������E��}� t\�}� tV�E�P�M誜���}� t=�E쉅������������������ tj�������n���� ����
ǅ ���    �E�    �E�R��P���Kr��XZ_^[��   ;�蓆����]� �   �����   �str ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P��q�����E�_^[���   ;��څ����]� ������������������������U���  SVWQ�������B   ������Y�M��M������E�P�MQ�M�輚���Eԃ}� uǅ����    �M������������#�E�P�M�m���Eԉ�����M�还�������R��P�H��p��XZ_^[��  ;�������]�    P����   \str ������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��;�M�������P�EP�MQ�M�X{��P�U��BP��*�Q0�B<�Ѓ�;��a���_^[���   ;��Q�����]� �����������������������������������������������U����   SVWQ������9   ������Y�M��E�    �E�P�MQ�M���n���E��E�P�MQ�M�y���E�R��P���co��XZ_^[���   ;�諃����]� �   �����   �b ��������������������������������������������������U����   SVWQ������9   ������Y�M��E�P�MQ�M�輐���E��E�P�MQ�M�~���E�R��P�p�n��XZ_^[���   ;�������]�    x����   �b ������������������������������������������U����   SVWQ������:   ������Y�M��E�P�MQ�M������E܃��E��$�EP�M�i���E�R��P�(��m��XZ_^[���   ;��=�����]� �I    0����   <b ��������������������������������������������������U����   SVWQ������;   ������Y�M��M�������E�P�MQ�M��'�����u3��E�E�P�MQ�M�������u3��-�E�P�MQ�M��������u3���E�P�MQ�M��r���   R��P� ��l��XZ_^[���   ;��C�����]� �   (����   4v ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E����X�M����Y�U�����E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��PH��;��G���_^[���   ;��7�����]� �������������������������������������U����   SVWQ������?   ������Y�M��M��b����E�P�MQ�M������EԍE�P�MQ�M�ɒ���Eԉ�����M��+��������R��P���>k��XZ_^[���   ;������]�    �����   �b ����������������������������������������������U���  SVWQ�������B   ������Y�M��M�蚇���E�P�MQ�M��7����EȍE�P�MQ�M�x���Eȉ������M��6l��������R��P���nj��XZ_^[��  ;��~����]�    �����   �b ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P<��;��'~��_^[���   ;��~����]� �������������������������������������U���  SVWQ�������B   ������Y�M��M�������E�P�M�Q�UR�M���s���E��}�t�E�P�MQ�M��n���}�t���E��$�EP�M�d���E�R��P��i��XZ_^[��  ;��U}����]� �I    ����   2����   0b c ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�j j �EP�M��v��P�MQ�M��n��_^[���   ;��|����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��4|��_^[���   ;��$|����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E$P�M Qj �UR�EP�MQj �UR�M�x��P�EP�M��-���_^[���   ;��{����]�  ��������������������������������������U����   SVWQ��4����3   ������Y�M�j �E@P���E8�$���E0�$�M,Q���E$�$���E�$���E�$�����$�UR�M�it�����$�EP�M��}l��_^[���   ;���z����]�< ������������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP��*�Q�M����   ��;��_z��_^[���   ;��Oz����]� �����������������������������U����   SVWQ��4����3   ������Y�M�j ���E$�$���E�$���E�$�����$�EP�M�Cs�����$�MQ�M���m��_^[���   ;��y����]�$ ������������������������������������U����   SVWQ��4����3   ������Y�M�j ���E$�$���E�$���E�$�����$�EP�M�r�����$�MQ�M�����_^[���   ;��y����]�$ ������������������������������������U����   SVWQ��4����3   ������Y�M�j ���E$�$���E�$���E�$�����$�EP�M�r�����$�MQ�M���m��_^[���   ;��vx����]�$ ������������������������������������U���  SVWQ�������B   ������Y�M��EPj ������~��P�MQ�� ���R�M����P�EP�M��)s���������� ����d���������Y���������_^[��  ;���w����]� �����������������������������������U���   SVWQ�������H   ������Y�M�j ����������P�EP�����Q�M�rg��P�UR�M���z��������������d���������d��������_^[��   ;��w����]� ���������������������������������������U����   SVWQ������<   ������Y�M���EP�MQ�����R��*�P�M����   ��;��v��P�M腁���������c���E_^[���   ;��wv����]� �������������������������������������U���  SVWQ�������G   ������Y�M����]�}�t�����$�EP�M�uo���]�E P���E�$���E��$�������$y��P�MQ�����R�M�t[��P�EP�M������_^[��  ;��u����]� ���������������������������������������������������U����   SVWQ������;   ������Y�M���EP�MQ�����R��*�P�M����   ��;��.u���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;���t����]� ������������������������������������U���   SVWQ�������H   ������Y�M��} u��*�H�􋑘   ��;��t���E�} u3��  �M��f���E�htlfv�M��2c���M�i���M���$��a�����Mݝ�����k�����$��a����ܽ�������$hulav�M��7[��hmrffhtmrf�M��o���M�-i���M���$�a�����Mݝ�����Hk�����$�ta����ܽ�������$hinim�M���Z���M��h���M���$�Ba�����Mݝ������j�����$�&a����ܽ�������$hixam�M��Z�������$hpets�M��tZ��j hdauq�M��Gn���E�Phspff�M��6n���E Phsirt�M��%n���E�P�MQ������R�M��^�����\����������������}���M���[��������R��P��)�z^��XZ_^[��   ;���r����]�    �)����   �)msg ��������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U���  SVWQ�������C   ������Y�M��} u��*�H�􋑘   ��;��Jq���E�} u3��c�M�c���E�E�P�MQ�M�蘂���E��E��h���$�E��h���$�������:s���M���P�Q�P�Q�@�A�E�R��P��+�q\��XZ_^[��  ;��p����]� �I    �+����   �+b ��������������������������������������������������������������U����   SVWQ������?   ������Y�M�j �E P�MQ�UR������u��P�EP�� ���Q�M�Bv��P�UR�EP�M��^��_^[���   ;���o����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E�����E����X�E�_^[��]���������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R��*�P�M����   ��;��o���M���P�Q�P�Q�@�A�E_^[���   ;���n����]� ��������������������������������U����   SVWQ������<   ������Y�M��M��
t���E�P�MQ�UR�M��ox���EԍE�P�MQ�M�]���E�R��P�.�Z��XZ_^[���   ;��Vn����]�    .����    .time �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��P@��;���m��_^[���   ;��m����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��D�M�k����Pj j j j j j �M�d��Pj1�E��HQ��*�B0���   �у�(;��m��_^[���   ;��m����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj�E��HQ��*�B0���   �у�(;��cl���E�R��P�$0��W��XZ_^[���   ;��?l����]� �   ,0����   80r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��7��j j j j j j j �EPj-�M��QR��*�H0���   �҃�(;��k��_^[���   ;��uk����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��F�E�    ��E�Pj j j �MQ�URj j j)�E��HQ��*�B0���   �у�(;���j���E�R��P��1�mV��XZ_^[���   ;��j����]� �I    �1����   �1r ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��F�E�    ��E�Pj j �MQj �URj j j)�E��HQ��*�B0���   �у�(;���i���E�R��P��2�}U��XZ_^[���   ;���i����]� �I    �2����   �2r ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��=��j j j �EP�MQ�URj �EPj/�M��QR��*�H0���   �҃�(;���h��_^[���   ;���h����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj'�E��HQ��*�B0���   �у�(;��Ch���E�R��P�D4��S��XZ_^[���   ;��h����]� �   L4����   X4r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj,�E��HQ��*�B0���   �у�(;��Sg���E�R��P�45��R��XZ_^[���   ;��/g����]� �   <5����   H5r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj j �MQ�UR�EP�MQ�URj�E��HQ��*�B0���   �у�(;��cf���E�R��P�$6��Q��XZ_^[���   ;��?f����]� �   ,6����   86r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��M�E�    ��E�Pj �MQ�UR�EP�MQ�UR�EPj�M��QR��*�H0���   �҃�(;��re���E�R��P�7�Q��XZ_^[���   ;��Ne����]�    7����   (7r ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j �EP�MQ�URj �EPj.�M��QR��*�H0���   �҃�(;��d��_^[���   ;��d����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��*�B0���   �у�(;���c���E�R��P��8�wO��XZ_^[���   ;��c����]� �   �8����   �8r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj:�E��HQ��*�B0���   �у�(;���b���E�R��P��9�N��XZ_^[���   ;���b����]� �   �9����   �9r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��*�B0���   �у�(;��b���E�R��P��:�M��XZ_^[���   ;���a����]� �   �:����   �:r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj*�E��HQ��*�B0���   �у�(;��a���E�R��P�t;�L��XZ_^[���   ;���`����]� �   |;����   �;r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��*�Q0���   �Ѓ�(;��%`���E�R��P�d<�K��XZ_^[���   ;��`����]� �I    l<����   x<r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��*�Q0���   �Ѓ�(;��5_���E�R��P�T=��J��XZ_^[���   ;��_����]� �I    \=����   h=r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj	�U��BP��*�Q0���   �Ѓ�(;��E^���E�R��P�D>��I��XZ_^[���   ;��!^����]� �I    L>����   X>r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj
�U��BP��*�Q0���   �Ѓ�(;��U]���E�R��P�4?��H��XZ_^[���   ;��1]����]� �I    <?����   H?r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��*�B0���   �у�(;��c\���E�R��P�$@��G��XZ_^[���   ;��?\����]� �   ,@����   8@r ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��*�B0���   �у�(;��s[���E�R��P�A�G��XZ_^[���   ;��O[����]� �   A����   (Ar ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��=��j j j �EP�MQ�URj �EPj�M��QR��*�H0���   �҃�(;��Z��_^[���   ;��Z����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj�E��HQ��*�B0���   �у�(;���Y���E�R��P��B�gE��XZ_^[���   ;��Y����]� �   �B����   �Br ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��L�E�    ��E�Pj �MQ�UR�EP�MQj �URj>�E��HQ��*�B0���   �у�(;���X���E�R��P��C�wD��XZ_^[���   ;��X����]� �   �C����   �Cr ������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��*�Q0���   �Ѓ�(;���W���E�R��P��D�C��XZ_^[���   ;���W����]� �I    �D����   �Dr ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��H�M�U����Pj j j j �EP�MQ�M� N��Pj�U��BP��*�Q0���   �Ѓ�(;��W��_^[���   ;���V����]� ��������������������������������������������������U����   SVWQ������=   ������Y�M��EP�M���E���E�P�M�Q�M���V����t+�}� u��M��Pj��P�E�P�MQ�M��^����u3�����   R��P�<F��A��XZ_^[���   ;��(V����]� ��   DF����   pF����   lF����   hFdat sid br �������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��D�M��S����Pj j j j j j �M�4L��Pj�E��HQ��*�B0���   �у�(;��8U��_^[���   ;��(U����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E��x u3��J�E�    ��E�Pj j �MQ�UR�EPj �MQj�U��BP��*�Q0���   �Ѓ�(;��T���E�R��P�H�@��XZ_^[���   ;��aT����]� �I    H����   Hr ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��-��EP�MQ�UR�E��HQ��*�B0�HD�у�;��S��_^[���   ;��S����]� �����������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��EP�MQ�UR�EP�MQ�UR�E��HQ��*�B0�HH�у�;��S��_^[���   ;��S����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ��*�B0�HX�у�;��R��_^[���   ;��{R����]����������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)��EP�MQ�U��BP��*�Q0�BL�Ѓ�;��R��_^[���   ;���Q����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��)�E   ���P�M��QR��*�H0�QP�҃�;��sQ��_^[���   ;��cQ����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��$��EP�M��QR��*�H0�QP�҃�;���P��_^[���   ;���P����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��0��EP�MQ�UR�EP�M��QR��*�H0�QT�҃�;��LP��_^[���   ;��<P����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�HQ��*�B4��у�;���O���E�@    �E�M��H�M�
N����P�EP�MQ�M�rF��P�U��BP��*�Q0���   �Ѓ�;��xO���M�A�E3Ƀx ����_^[���   ;��TO����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��7��j j j j j �EPj j j�M��QR��*�H0���   �҃�(;��N��_^[���   ;��N����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��=�E�@    �M�QI����P�EP�M��BI��P��*�Q0���   �Ѓ�;��N��_^[���   ;��N����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j0�M��H��P��*�H0���   �҃�(;��M��_^[���   ;��rM����]�����������������������������������U����   SVWQ��4����3   ������Y�M��} u�E�*��EP�M�3��P�MQ�U��BP��*�Q0�B@�Ѓ�;���L��_^[���   ;���L����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��*�Q0�Bd�Ѓ�;��TL��_^[���   ;��DL����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��*�Q0�Bp�Ѓ�;���K��_^[���   ;��K����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��M�I����P�EP�MQ�UR�EP�M�B��P�M��QR��*�H0�Qh�҃�;��'K��_^[���   ;��K����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �M�A��Pj�E��HQ��*�B0���   �у�(;��J��_^[���   ;��|J����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j jj �M��@��Pj�E��HQ��*�B0���   �у�(;���I��_^[���   ;���I����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �M�H@��Pj�E��HQ��*�B0���   �у�(;��LI��_^[���   ;��<I����]� ������������������������������������������U���   SVWQ�� ����@   ������Y�M��M��K/���M�5G����P�E�Pj j j j j �M�?��Pj8�M��QR��*�H0���   �҃�(;��H���EЃ}� t�E�P�M��8���EЉ�����M��j1�������R��P�T�4��XZ_^[��   ;��OH����]� �   T����   (Tstorehere ��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�F����P�EPj j j j j �M�>��Pj9�M��QR��*�H0���   �҃�(;��G��_^[���   ;��tG����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��M�}E����Pj j j j j j �M��=��Pj"�E��HQ��*�B0���   �у�(;���F��_^[���   ;���F����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M��D����Pj j j j j j �M�A=��Pj5�E��HQ��*�B0���   �у�(;��EF��_^[���   ;��5F����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M�=D����Pj j j j �EPj �M�<��Pj<�M��QR��*�H0���   �҃�(;��E��_^[���   ;��E����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j j �EP�MQ�UR�EPj �MQj3�U��BP��*�Q0���   �Ѓ�(;��	E��_^[���   ;���D����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j �EPj �MQj�U��BP��*�Q0���   �Ѓ�(;��oD����EP�M��QR��*�H0�Qt�҃�;��KD��_^[���   ;��;D����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j �EPj j�M��QR��*�H0���   �҃�(;��C��_^[���   ;��C����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j�E��HQ��*�B0���   �у�(;��#C��_^[���   ;��C����]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j �EPj�M��QR��*�H0���   �҃�(;��B��_^[���   ;��B����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j(�E��HQ��*�B0���   �у�(;��B��_^[���   ;���A����]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j �EP�MQj&�U��BP��*�Q0���   �Ѓ�(;��oA��_^[���   ;��_A����]� �����������������������������U����   SVWQ��4����3   ������Y�M���j j j j �EP�MQj �URj+�E��HQ��*�B0���   �у�(;���@��_^[���   ;���@����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j�E��HQ��*�B0���   �у�(;��C@��_^[���   ;��3@����]������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j#�E��HQ��*�B0���   �у�(;��?��_^[���   ;��?����]������������������������������������U����   SVWQ��4����3   ������Y�M��} tj j�M�,<���M��} tj j�M�<���M���EP�MQ�U��BP��*�Q0�B`�Ѓ�;��?��_^[���   ;���>����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��*�B0���   �у�;��i>��_^[���   ;��Y>����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j �E��HQ��*�B0���   �у�(;���=��_^[���   ;���=����]������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��M��<���E�� x�E��@   �E��@    �E�_^[���   ;��;����]����������������������������������U����   SVWQ��4����3   ������Y�M��M���4���E��t�E�P�'�����E�_^[���   ;��
;����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� x�M��79��_^[���   ;��:����]�������������������������U����   SVWQ��0����4   ������Y�M��E��@    j �EP�MQ�UR�EPj 3Ƀ} ����
Q�M������t�U��z tǅ0���   �
ǅ0���    ��0���_^[���   ;���9����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�M��<��_^[���   ;��9����]� ����������������������U����   SVWQ������:   ������Y�M��M�l'������������ckhc)�����ckhct5�����cksatY�����TCAbtr��   �����atnit��   3���   �E��x t �M��9����t�E��@    �   �   3��   �E��x t�E����M��B��;��8���}3��yj hdiem�M�o5���E�E��@   ��EP�M�Q�U���M��P��;��_8���E��E��x t�}�t�}�u3��}���P�M��F���E���EP�MQ�M��,��_^[���   ;��8����]� ����������������������������������������������������������������������������������������������U����   SVWQ�� ����8   ������Y�M��E��x u�  �E�� ����� �����   �� ����$� f�E;E~��   �   �E;E|��   �{�E;E}�   �l�E;E�   �]�E;E~�E;E}�   �F�E;E|
�E;E�|�2�E;E|
�E;E}�h��E;E~
�E;E�T�
�E;Et�H�EP��(����6����(���Q�M��29��j�E���$�E���$�EP��K�����E��@    _^[���   ;��d6����]� ��ee%e4eCeZene�e�e������������������������������������������������������������������������������������������������������������U����   SVWQ�� ����8   ������Y�M��E��x u�X  �E�� ����� �����   �� ����$�0h�E�]����z�#  ��   �E�]����Az�  �   �E�]����Au��   �   �E�]����u��   �   �E�]����z�E �]����Au�   �n�E�]����Az�E �]����u�   �M�E�]����Az�E �]����Au�{�/�E�]����z�E �]����u�]��E�E������D{�J�EP��(����y4����(���Q�M��7���E(P���E �$���E�$�MQ�I�����E��@    _^[���   ;��34����]�$ ��f�fg)g@gag�g�g�g����������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�j���E �$���E�$���E�$�EP�MQ�M�����_^[���   ;��,3����]�  ��������������������������U����   SVWQ��4����3   ������Y�M�j���E �$���E�$���E�$�EP�MQ�M��Y��_^[���   ;��2����]�  ��������������������������U����   SVWQ��4����3   ������Y�M�j���E �$���E�$���E�$�EP�MQ�M�����_^[���   ;��,2����]�  ��������������������������U����   SVWQ��4����3   ������Y�M��E�� ��E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��l'���E��t�E�P�L�����E�_^[���   ;��J1����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� ��E��x u ��E��HQ��*�B4��у�;���0���E��@    �E��@    _^[���   ;��0����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Qt�҃�;��E0��_^[���   ;��50����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��} tT��EP�M���*��P��*�Q0���   �Ѓ�;��/���E��EP�M�Q��*�B0���   �у�;��/���$��EP�M��QR��*�H0�Q|�҃�;��k/��_^[���   ;��[/����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H�у�;���.��_^[���   ;���.����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H�у�;��h.��_^[���   ;��X.����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H�у�;���-��_^[���   ;���-����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H|�у�;��-��_^[���   ;��x-����]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4���   �у�;��-��_^[���   ;��-����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4�Q�҃�;��,��_^[���   ;��y,����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4�Q�҃�;���+��_^[���   ;���+����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�Q/����u�M���P�M��<���6�M�1/����u�M�:��P�M��H���h�����P������_^[���   ;��3+����]� �������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �B@�Ѓ�;��*��_^[���   ;��*����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Q �҃�;��E*��_^[���   ;��5*����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Q$�҃�;���)��_^[���   ;��)����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H0���   �҃�;��6)��_^[���   ;��&)����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4���   �҃�;��(��_^[���   ;��(����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��*�Q4���   �Ѓ�;��!(��_^[���   ;��(����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��BP��*�Q4���   �Ѓ�;��'��_^[���   ;��'����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Q(�҃�;��'��_^[���   ;��'����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��*�B4�H,�у�;��&��_^[���   ;��|&����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�B0�Ѓ�;��&��_^[���   ;�� &����]� ������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H4�у�;��%��_^[���   ;��%����]�������������������������U���(  SVWQ�������J   ������Y�M��E�    �E�    �E�P�M�Q�UR�E��H��5���M���5��P�������%���E�P�M�Q�U�R�E�P������Q�U��J�58���} tL�} tF�E�;E�~*�M�M�9M�}�U�;U�~�E�E�9E�}ǅ����   �
ǅ����    �������h�7�} t1�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    �������/�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    ������R��P�Px����XZ_^[��(  ;��$����]� �I    Xx����   �x����   �x����   �x����   �x����   �x����   �xdy dx h w y x ������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Q8�҃�;���"��_^[���   ;���"����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Q<�҃�;��u"��_^[���   ;��e"����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4���   �Ѓ�;���!��_^[���   ;���!����]� ���������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H@�у�;��x!��_^[���   ;��h!����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�BD�Ѓ�;�� !��_^[���   ;��� ����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�BH�Ѓ�;�� ��_^[���   ;��p ����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�BL�Ѓ�;��  ��_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�BP�Ѓ�;����_^[���   ;��p����]� ������������������������������U����   SVWQ��4����3   ������Y�M��M��"������   �M��"����u5�M�����P�M���P�E��HQ��*�B4�HP�у�;������X�M�"����u5�M�.����P�M����P�E��HQ��*�B4�HH�у�;�����h�����P�4������   �M�1"������   �M� "����u5�M�j����P�M�-��P�E��HQ��*�B4�HL�у�;��(���X�M��!����u5�M�k-����P�M�`-��P�E��HQ��*�B4�HD�у�;������h�����P������h�����P�l����_^[���   ;������]� ��������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4��  �҃�;�����_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�M��QR��*�H4�QT�҃�,;��1��_^[���   ;��!����]�( �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4�QX�҃�;����_^[���   ;������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H`�у�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�Hd�у�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4��   �҃�;��&��_^[���   ;������]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E��HQ��*�B4�H\�у�;����_^[���   ;������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�Bh�Ѓ�;����_^[���   ;�� ����]� ������������������������������U����   SVWQ��(����6   ������Y�M��} t�E��ًU�
�} t�E��ًU�
��EP�MQ�U��BP��*�Q4�Bh�Ѓ�;��l���E�} t�E��ًU�
�} t�E��ًU�
�E�_^[���   ;��2����]� ������������������������������������������������U����   SVWQ��(����6   ������Y�M��} t�E��ًU�
�} t�E��ًU�
��EP�MQ�U��BP��*�Q4�Bp�Ѓ�;�����E�} t�E��ًU�
�} t�E��ًU�
�E�_^[���   ;��R����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�Bp�Ѓ�;�����_^[���   ;�������]� ������������������������������U���  SVWQ�������D   ������Y�M��E��x ��   �} t1�M��'����P�E��H�d��P��*�Q0�Bl�Ѓ�;��7���T�M���&��P��������hARDb����������P�����P�� ���Q�U��J�p���� ���� �������������_^[��  ;�������]� ���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR��*�H4�Ql�҃�;��E���   _^[���   ;��0����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$���E�$�MQ�U��BP��*�Q4���   �Ѓ�;����_^[���   ;������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��*�B4���   �у�;����_^[���   ;��	����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4���   �у�;����_^[���   ;������]��������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M�h�  �M�����EP�MQ�UR�EP�M��5!��2�_^[���   ;������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M���M��B��;����_^[���   ;������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR��*�H4�Qx�҃�;��I��_^[���   ;��9����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�UR�E��H����_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M��} tj j�M�L���M��} tj j�M�5���M���EP�MQ�U��BP��*�Q4�Bp�Ѓ�;��"��_^[���   ;������]� ������������������������������������������������U���0  SVWQ�������L   ������Y�M��E�    �M�����������������INIbf������INIb��   ������SACb5������SACb��   ������$'  ��  ������MicM��  �$  ������ARDb�4  �  ������NIVb1������NIVbt\������NPIb�v  ������ISIb��   ��  ������cnys��  �  �E����M��B��;������E�   �  �E����M��B��;�����E�   �y  �E�    �E�    ��E�P�M�Q�U���M��P��;��p����t)��E�P�M�Q�U��BP��*�Q4�B�Ѓ�;��C���E�   �  �M�������P�M�����P�E���M��B��;�����E�   ��   j j�M��	���E�j j�M��	���E�j j�M�	���E�j j�M�	���E���EP�M�Q�U�R�E�P�M�Q�U���M��P��;�����E�   �q��EP�M���M��B��;��z���X��EP�M���M��B$��;��^���E�   �2j hIicM�M�+	���E��EP�M�Q�U���M��P ��;��%����E�R��P�d�����XZ_^[��0  ;�������]� �   l�����   ������   ��h w ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�h����h����h�����EP�MQh����h����h����h�����UR�M������_^[���   ;��
����]� ��������������������������������U����   SVWQ������:   ������Y�M�hYALf���������P�M�����������)���_^[���   ;��%
����]��������������������������������������U����   SVWQ��4����3   ������Y�M��M���
���E�� 0�E��@   �E�_^[���   ;��	����]����������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�<������E�_^[���   ;��:	����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� 0�M��g��_^[���   ;�������]�������������������������U����   SVWQ��0����4   ������Y�M��M������0�����0���cksat9��0���ckhct�P�E��@   �M������t�E��@    �   �93��5�E��x t�E����M��B��;��'���3���EP�MQ�M��	���_^[���   ;������]� ���������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��*�H���  �҃�;��j��_^[���   ;��Z����]���������������������������U����   SVW��@����0   �������EP��*�Q0���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��(����6   �������EP�MQ��,���R��*�H0���   �҃�;����P�M������,��������E_^[���   ;��\����]���������������������������������������������U���,  SVW�������K   ������M�����E�    �	�E����E�   ����   j �E�k�
P�M����E�j �E�k�
��P�M����Eȃ}� u�b�}� ~,j h\���������������P�M����������� ���E�P�M�Q������R�?����P�M��Y�������������U����E�P�M�����M�����ER��P�H������XZ_^[��,  ;������]Ë�   P�����   \�t ����������������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ��*�B0���   �у�;��i��_^[���   ;��Y����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR��*�H0���   �҃�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   ������j0j �b����P�EP�����_^[���   ;��u����]����������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVW��@����0   ������j0j ������P�EP������P�b����_^[���   ;�������]�����������������������������U����   SVW��(����6   ������j0j �R����P�EP�MQ��,���R�k�����P��������,�������_^[���   ;��F����]���������������������������������������U����   SVW��(����6   ������j0j ������P�EP�MQ�UR��,���P������P�S������,����@��_^[���   ;������]�����������������������������������U����   SVW��@����0   ������j j�2����P�EP������3Ƀ�����_^[���   ;��;����]����������������������������U����   SVW��@����0   ������j j������P�EP������P�b����3Ƀ�����_^[���   ;��� ����]�����������������������������������U����   SVW������9   ������j j�B����P�EP�MQ��,���R�[�����P������3Ƀ����� �����,�������� ���_^[���   ;��" ����]�����������������������������������U����   SVW������9   ������j j�
����P�EP�MQ�UR��,���P�������P�3����3Ƀ����� �����,�������� ���_^[���   ;��~�����]�����������������������������������������������U����   SVW��@����0   �������EP�MQj ��*�B���   �у�;�����_^[���   ;��������]������������������������U����   SVW��@����0   �������EP�MQ�URj ��*�H���   �҃�;�����_^[���   ;�������]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E��HQ��*�B4�H,�у�;�����_^[���   ;��������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��BP��*�Q4�B0�Ѓ�;�����_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�B4�H4�у�;�����_^[���   ;�������]�������������������������U����   SVWQ������9   ������Y�M��M����� �E�M�����E��}� t�E�   �E�P�M�Q�UR�M�����_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M��E P�MQ�M����P�UR�EP�MQ�M�����R�EP�M����_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��M����P�E<P���E4�$���E,�$�M(Q���E �$���E�$���E�$�M�������� �$�UR�M������_^[���   ;��?�����]�8 ���������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����P���E �$���E�$���E�$�M�H������ �$�EP�M�����_^[���   ;�������]�  ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�4���P���E �$���E�$���E�$�M������� �$�EP�M�����_^[���   ;��������]�  ���������������������������������������U����   SVWQ��4����3   ������Y�M��M����P���E �$���E�$���E�$�M������� �$�EP�M�����_^[���   ;��Y�����]�  ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�����P�EP�MQ�UR�M�X���P�EP�MQ�M��o���_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M��EP�M�r���P�M����P�MQ�M�����_^[���   ;��W�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E P���E�$���E�$�M�����P�MQ�M����_^[���   ;��������]� ����������������������������U���  SVWQ�������F   ������Y�M��E�P�M�Q�UR�M��#���E�P�M�Q�U�R�E�P�MQ�M��
���} tL�} tF�E�;E�~*�M�M�9M�}�U�;U�~�E�E�9E�}ǅ����   �
ǅ����    �������h�7�} t1�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    �������/�E�;E�~�M�M�9M�}ǅ����   �
ǅ����    ������R��P���8���XZ_^[��  ;�������]� ��   �����   @�����   >�����   <�����   :�����   7�����   4�dy dx h w y x ��������������������������������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E�E�}� u	�E����E�j hdiuM�M�J����E��}� u�   �G�E�M�;u3��9j hIicM�M����9E�uj h1icM�M������t3���E�M���   _^[���   ;��������]� ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M����   ��;��t���_^[���   ;��d�����]� ����������������������������������U����   SVW������:   ������hfnic�M�Q����E��}� tj
�M�������t�\hfnic�����P�M�����P�M�@��������������M��������t�M�������uhfnic�M������EPj
�M���_^[���   ;�������]�������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��B$��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ������:   ������Y�M���EP�����Q��*�B�M��PP��;��$���P�M��������������E_^[���   ;��������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�M��BT��;�����_^[���   ;��{�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��3���P��*�Q0���   �Ѓ�;�����_^[���   ;��������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M�������Pj j j �EP�MQj �M�]���Pj=�U��BP��*�Q0���   �Ѓ�(;��a���_^[���   ;��Q�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��M�M�����P�EPj j j��MQj �M����Pj=�U��BP��*�Q0���   �Ѓ�(;�����_^[���   ;�������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���j j j j j j j j j6�M��A���P��*�H0���   �҃�(;�����_^[���   ;�������]�����������������������������������U����   SVWQ��(����6   ������Y�M�j �EP�M������E�E�P�M��$���_^[���   ;�������]� ��������������������������U����   SVWQ��(����6   ������Y�M�j �EP�M� ����E�E�P�M������_^[���   ;�������]� ��������������������������U����   SVWQ��$����7   ������Y�M������$�EP�M�0����]���E��$�M�����_^[���   ;�������]� �������������������������������U���,  SVWQ�������K   ������Y�M��M���������������P�EP������Q�M�������U؋H�M܋P�U��H�M�P�U�@�E���ċM؉�U܉P�M��H�U�P�M�H�U�P�M��T���R��P����v���XZ_^[��,  ;�������]�    ������   ��val ��������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M���������������P�EP�����Q�M�H�����U��H�M�P�U�@�E���ċM���U�P�M�H�U�P�M������R��P����n���XZ_^[��  ;�������]�    ������   ��val ������������������������������������������������������������U���   SVWQ�������H   ������Y�M��M���������������P�EP������Q�M����P�M�� ���������|����������q������̍E�P�g����M�������M��S���R��P����l���XZ_^[��   ;�������]� ��   ������   ıval ��������������������������������������������������������U����   SVWQ������:   ������Y�M��E;Eu&j htsem�M������uj hrdem�M�������t3��B�E�    �EP�����������M�Q�����R�M�������u3���E�P�M��R����   R��P����\���XZ_^[���   ;�������]� ��   Ȳ����   Բval ��������������������������������������������������������U����   SVWQ������:   ������Y�M��E;Eu&j htsem�M�������uj hrdem�M�������t3��B�E�    �EP�����������M�Q�����R�M�a�����u3���E�P�M��c����   R��P�г�L���XZ_^[���   ;�������]� ��   س����   �val ��������������������������������������������������������U����   SVWQ������;   ������Y�M��E;Eu&j htsem�M�������uj hrdem�M�������t3��E���]�EP�����������M�Q�����R�M�6�����u3�����E��$�M������   R��P���9���XZ_^[���   ;�������]� �I    �����   ��val ��������������������������������������������������������������������U���  SVWQ�������G   ������Y�M��E;Et�E;Et�E;Et3���   j htsem�M������uj hrdem�M������t3��   �����$�M������EP�����������MQ�������z����UR������k����E�P������Q������R�����P�M�������u3��5���ċM؉�U܉P�M��H�U�P�M�H�U�P�M������   R��P�t�����XZ_^[��  ;��������]� �I    |�����   ��val ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X�M��E�Y�U��E��E�_^[��]� �����������������������U����   SVWQ������=   ������Y�M��E;Eu&j htsem�M�������uj hrdem�M������t3��_�M��(����EP����������M�Q�UR�����P�M�{�����u3��)���ċM���U�P�M�H�U�P�M������   R��P�������XZ_^[���   ;��G�����]� �   $�����   0�val ����������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��E;Eu&j htsem�M������uj hrdem�M�t�����t3��v�M�� ����EP�������k����M�Q������R�M������uǅ����    �M�������������.���̍E�P�����M��7���ǅ���   �M����������R��P�t�����XZ_^[��  ;��������]� ��   |�����   ��val ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������E�� d�E��M�Hj hmyal�M�%����M��A�E��xt�E��xt
�E��@    j
hhfed�M������M��A�E�_^[���   ;��������]� ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�l������E�_^[���   ;��j�����]� ������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;�������]������������������U����   SVWQ��0����4   ������Y�M��M�������0�����0���ytsdt�%�M�������E����M��B��;������   ��EP�MQ�M�����_^[���   ;��x�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ������;   ������Y�M��M�������E�P�M�#����M��b����ER��P�<������XZ_^[���   ;��)�����]� �I    D�����   P�tri ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M����l���_^[���   ;�������]�������������������������������U����   SVWQ��4����3   ������Y�M��E��M���E��P�M��������E�_^[���   ;��*�����]� ������������������������U����   SVWQ��4����3   ������Y�M��E����M��BD��;��������t*�E��H;Mt�E��M�H�E����M��BH��;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��x u3���E��H��������_^[��]�������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M���_^[��]������������������U����   SVWQ��4����3   ������Y�M������$�E��H������E�P�M��Q�E��H��B$��;������j j h����(�����_^[���   ;��������]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X(_^[��]� ���������������������������U���l  SVWQ�������[   ������Y�M��􍅘���P�M���M��B(��;�����P�M��0�������������j �������|���Pj jj?j �M�������������]���j �������S���Pj j(������Pjh�  �M��}��������������������������������t3���   j �����������Pj j j8j �M����������������j�M��,��������跿��Pj�;�����Ph,  �-�����Pj;�� �������Ph	��h�  �M��~����� ������������������M��1����M��)���j�M��j����E��M��H$j�������   _^[��l  ;�������]������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������j �EP������_^[���   ;�������]�����������������U����   SVW��@����0   ������E��E_^[��]�������������������U����   SVWQ������=   ������Y�M�j�M����*����E��@4    �E��@8    �E��@<    �E����X(h�   �M�����j h�������V���h�  ��(����2���j j �����P��(���Q�M��O������������j j�M��������_^[���   ;��������]����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��(����6   ������Y�M��E�    �   ����   �E��x4 t8h��0��P�ܾ����j
�+������M����*�����t3��   뿋M���0������E��x4 ur�E��M�H8�E��M�H4�M���0������E��x4 tj
��������M����������t3��X�؋M���0�����E��H<�M�E��@<    �M���0�{����(�!h��0��$P�������M���0�V��������E�_^[���   ;��E�����]� �����������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���*�PP��M��Bh��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���*�PP��M��Bl��;��@���_^[���   ;��0�����]���������������������������������U����   SVWQ��4����3   ������Y�M���E��HQ��*�BP�H�у�;������_^[���   ;�������]�������������������������U���h  SVWQ�������Z   ������Y�M�j h��������v���h�  �������R���j j ������P�M��A(�X����P������R�b�����P������P�!�����P������Q�M��=����������~����������s����������h���htats�M�����jj�M��	����E����@(�$j�M��޹��h�  �����������E�P������Q�����R�M��
���������D����E��x4 tl�M���0�a����E��x4 t7��E��H8Q�U��B4�Ѓ�;��N����M��A<�E��@8    �E��@4    �h��4��P�Һ�����M���0�
����M������R��P�|�蠽��XZ_^[��h  ;��������]� ��   ������   ��m ������������������������������������������������������������������������������������������������������������������������������U���0  SVWQ�������L   ������Y�M��M�L���������������MicMtM������fnict�   j�����������P�M�M����������ѹ��jj�M������   �   �   j hIicM�M�������������������t�`htats�M��b���j j�M�����h�  �������q����E�P������Q�����R�M��ջ������������M��=���j�M������EP�MQ�M��r���R��P�T��ƻ��XZ_^[��0  ;�������]�    \�����   h�m ��������������������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��0�����0���t�(j�M��������j�,�����j �M������   ��EP�MQ�M�覿��_^[���   ;�������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M�j�M����Z���j������3�_^[���   ;�������]���������������������������������U����   SVWQ������9   ������Y�M��M���賴���E�� ������ ���蟴��P�M����u����� ���������E�_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M�j �E�P�M�����E�_^[���   ;��X�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�UR��*���   �Q�҃�;������_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �EP�M��������$�E��8 u�EP�M����������t	�E��    �M�)���_^[���   ;�������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����������_^[���   ;��'�����]� ���������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u�E��     �E��E�X�#�E��8 u�E��@�E������D{	�E��    _^[��]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u4�E��     �E����M��U�P�M�H�U�P�M�H�U�P�(�E��8 u �EP�M���Q�۬������t	�E��    _^[���   ;�������]� ���������������������������������������������������U����   SVW��<����1   ������E�M� �������Dz6�U�E�B�@������Dz!�M�U�A�B������Dzǅ<���    �
ǅ<���   ��<���_^[��]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�3Ƀ8����_^[��]��������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8�u(�E��     �E����M��U�P�M�H�U�P�(�E��8 u �EP�M���Q��������t	�E��    _^[���   ;�������]� �����������������������������������������������U����   SVW��4����3   ������E�M� �������Dz�E�M�@�A������Dz3��c�E�M� �I���$� ������U�E��H���$ݝ8���������݅8���������D{ǅ4���   �
ǅ4���    ��4���_^[���   ;�������]����������������������������������������������������������������U����   SVW��@����0   ������E�8 t��E�Q��*�B��у�;������E�     _^[���   ;��~�����]�������������������������������U����   SVW��@����0   �������hﾭޡ�*�H��@  �҃�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   ������} t!��EP��*�Q��@  �Ѓ�;�����_^[���   ;�������]������������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;��9���_^[���   ;��)�����]��������������������������U����   SVW��@����0   �������EP�MQ��*�B��  �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �����󫡘*�H��   ��;��e���_^[���   ;��U�����]����������������������U����   SVW��@����0   ������} t�E�x��u�   �3�_^[��]��������������������U����   SVW��<����1   ������=�* tE�}sǅ<���   �	�E��<�����j j ��<���Q��*�B���   �у�;������j�EP�I   ��_^[���   ;��b�����]���������������������������������������������������U����   SVW��4����3   ������}s�E   �E��P�/������E��}� u3��:�} t�E��Pj �M�Q��������E�� �����E����E���*   �E�_^[���   ;�蛿����]��������������������������������������������U����   SVW��<����1   ������=�* tE�}sǅ<���   �	�E��<�����j j ��<���Q��*�B���   �у�;������j�EP�������_^[���   ;�������]���������������������������������������������������U����   SVW��<����1   ������=�* tE�}sǅ<���   �	�E��<�����j j ��<���Q��*�B���   �у�;��B����j�EP�	�����_^[���   ;��"�����]���������������������������������������������������U����   SVW��<����1   ������=�* tE�}sǅ<���   �	�E��<�����j j ��<���Q��*�B���   �у�;�肽���j�EP�I�����_^[���   ;��b�����]���������������������������������������������������U����   SVW��4����3   ������} tF�E�E��=�* t�E�x��u�E��P���������E�P��*�Q��Ѓ�;��¼��_^[���   ;�貼����]�����������������������������������U����   SVW��4����3   ������} tF�E�E��=�* t�E�x��u�E��P�e��������E�P��*�Q��Ѓ�;��"���_^[���   ;�������]�����������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;�豻��_^[���   ;�衻����]����������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;��A���_^[���   ;��1�����]����������������������������������U����   SVW��<����1   ������=�* tI�}sǅ<���   �	�E��<�����MQ�UR��<���P��*�Q���   �Ѓ�;�螺���j�EP�e�����_^[���   ;��~�����]�����������������������������������������������U����   SVW��<����1   ������=�* ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P��*�Q���   �Ѓ�;��Թ���[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P��*�Q���  �Ѓ�;�艹����EP�MQ�N�����_^[���   ;��g�����]������������������������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�* t0��EP�MQ�UR��*�H���   �҃�;��������0����j�EP��������0�����0����M��E���th��8��
P�3������E�_^[���   ;��j�����]�����������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�* to�} t0��EP�MQ�UR��*�H���   �҃�;��ʷ����0����.��EP�MQ�UR��*�H���  �҃�;�蚷����0�����0����E��j�EP�R������E��E���th��<��P�������E�_^[���   ;��G�����]������������������������������������������������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;������_^[���   ;�豶����]����������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;��Q���_^[���   ;��A�����]����������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;�����_^[���   ;��ѵ����]����������������������������������U����   SVW��@����0   �������EP��*�Q��Ѓ�;��q���_^[���   ;��a�����]����������������������������������U����   SVW��@����0   �������EP��*�Qp��Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������h   ��*�Hp��҃�;�葴��_^[���   ;�聴����]����������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��*�Bp�H�у�;������E�     _^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�Hp�Q�҃�;�蔳��_^[���   ;�脳����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�Hp�Q�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�Hp�Q�҃�;�蔲��_^[���   ;�脲����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�Bp�H�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �   ���E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��p���_^[���   ;��`�����]� ����������������������������������������������U����   SVW��@����0   ������h�*�EPhD �9�����_^[���   ;�������]�������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��d���_^[���   ;��T�����]� ����������������������������������U����   SVWQ������>   ������Y�M�h�   ��������E�}� t�E샸�    u3��?�M��]����E�P�MQ�e�������u3����EP�M�Q�U�M����   ��;�褯��R��P����;���XZ_^[���   ;�胯����]� �   ������   ��dat ��������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��Į��_^[���   ;�贮����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u���EP�U�M����   ��;��*���_^[���   ;�������]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u���EP�U�M����   ��;�芭��_^[���   ;��z�����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u���EP�U�M����   ��;�����_^[���   ;��ڬ����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u���EP�U�M����   ��;��J���_^[���   ;��:�����]� ����������������������������������������U����   SVWQ������9   ������Y�M���EP��*�Q�M��Bd��;��˫���E�}� u3��s��h8�@��P�M��Q��*�B���   �у�;�茫���E��}� u3��4��EP�M��Q�U�R��*�P�M��Bh��;��W����E�E��  �E�_^[���   ;��;�����]� ���������������������������������������������������������U����   SVW��@����0   ������j h�  h�*�M������*_^[���   ;�赪����]����������������������U����   SVW��@����0   ������j h�  h�*�M赯����*_^[���   ;��U�����]����������������������U����   SVW��@����0   ������h� �M貚����tj h�  h�*�M踚�����=����h�h�*�Ԙ������*_^[���   ;��ɩ����]������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M��B��;��X���_^[���   ;��H�����]� ����������������������U����   SVWQ��4����3   ������Y�M���*���   ��M��Bx��;�����_^[���   ;��ݨ����]������������������������������U����   SVW��(����6   ������j h�  h�*��,���P�M肐�����ǭ����,���������*_^[���   ;��\�����]�����������������������������U����   SVW��(����6   ������j h�  h�*��,���P�M�������G�����,����o�����*_^[���   ;��ܧ����]�����������������������������U���  SVW�������B   ������h3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |I�E�M������E��E���
}�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�먋E��D� j �E�P�M������ER��P���肒��XZ_^[�M�3��*�����  ;��������]�   ������   ��hexstring ����������������������������������������������������������������������������������U���  SVW��x����b   ������} ��   �}   @��   j h�����������Pj0j jj �E�U��m�����x�����|���߭x����5����$������P�]�����P�MQ蹶�����������&��������������E�^  �  �} ��   �}   ��   j h��������t���Pj0j jj �E�U�
�ώ����x�����|���߭x����5����$������P迺����P�MQ������������舸���������}����E��   �r�} |l	�}   vaj h�����������Pj0j jj �m�5����$������P�H�����P�MQ褵�������������������������E�Lj h������耮��P�EP��,���Q蔬����P�UR�V�������,����÷�������踷���E_^[�Ĉ  ;��'�����]��������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   ��������E P�MQ�UR�EP���E�$��,���Q��*�B�H$�у�;��3���P�M謭����,���蝶���E_^[���   ;�������]���������������������������������������������U����   SVW��4����3   ������j�   ���E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;��m���_^[���   ;��]�����]����������������������������������������������U����   SVW��@����0   ������hX/�EPh�f �9�����_^[���   ;�������]�������������������������U����   SVW������<   ������j�{������E��}� t	�E��x uǅ��������M�َ��������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�F����EP�M��Q�҃�4�� ����M蒎���� ���_^[���   ;��#�����]����������������������������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;�蒠��_^[���   ;�肠����]�����������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�M��Q�҃�;�����_^[���   ;��������]���������������������������������������U����   SVW��@����0   �����󫡘*�HL���   ��;�蕟��_^[���   ;�腟����]����������������������U����   SVW��@����0   �������E�Q��*�B@�H�у�;��.����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �����󫡘*�HL����;�蹞��_^[���   ;�詞����]��������������������������U����   SVW��@����0   �������E�Q��*�B@�H�у�;��N����E�     _^[���   ;��5�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL���   �Ѓ�;��ȝ��_^[���   ;�踝����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL���   �҃�;��Q���_^[���   ;��A�����]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P��*�QL���   �Ѓ�;��؜���E�}� u)��j �EP�M�Q��*�BL���   �у�;�訜����M������P�M觲��_^[���   ;�腜����]� ���������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M��BH��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���*���   ��M��BP��;�蝛��_^[���   ;�荛����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL��(  �Ѓ�;��(���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL��,  �҃�;�豚��_^[���   ;�衚����]� �������������������������������U����   SVW��@����0   �����󫡘*�HL��Q��;��H���_^[���   ;��8�����]�������������������������U����   SVW��@����0   �������E�Q��*�B@�H�у�;��ޙ���E�     _^[���   ;��ř����]��������������������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R��*�HL�Q�҃�;��Q���P�M�͖��������1����E_^[���   ;��*�����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL���   �у�;�贘��_^[���   ;�褘����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL�Q�҃�;��4���_^[���   ;��$�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B�Ѓ�;�軗��_^[���   ;�諗����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B�Ѓ�;��K���_^[���   ;��;�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B�Ѓ�;��ۖ��_^[���   ;��˖����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�QL�B �Ѓ�;��_���_^[���   ;��O�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL��4  �у�;�����_^[���   ;��ԕ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�QL�B$�Ѓ�;��_���_^[���   ;��O�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�BL�H(�у�;��۔��_^[���   ;��˔����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B,�Ѓ�;��k���_^[���   ;��[�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B0�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL��  �҃�;�聓��_^[���   ;��q�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL���   �Ѓ�;�����_^[���   ;��������]�������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R��*�HL��  �҃�;�莒��P�M�
���������n{���E_^[���   ;��g�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B4�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P��*�QL�B8�Ѓ�;�艑��_^[���   ;��y�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�蔐��_^[���   ;�脐����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�蔏��_^[���   ;�脏����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�BL�M����   ��;�蔎��_^[���   ;�脎����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�QL�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�QL�M����   ��;�訍��_^[���   ;�蘍����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�QL�M����   ��;��8���_^[���   ;��(�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL�H<�у�;��ǌ��_^[���   ;�跌����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B�Ѓ�;��K���_^[���   ;��;�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL�Q@�҃�;��ԋ��_^[���   ;��ċ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q��*�BL�HD�у�;��U���_^[���   ;��E�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q��*�BL�HH�у�;��Պ��_^[���   ;��Ŋ����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q��*�BL�HD�у�;��U���_^[���   ;��E�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q��*�BL�HH�у�;��Չ��_^[���   ;��ŉ����]� �����������������������������������U���,  SVWQ�������K   ������Y�M��M���o��h�  �������vy��P�������{��j �E�P������Q�M��hp��������������������N�����������tǅ���    �M��ɓ���������M��U���������M�諓�������R��P���~t��XZ_^[��,  ;��ƈ����]Ë�   �����   �dat ����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U���  SVWQ�������B   ������Y�M�j�������U���h�  ��$�����w��P������z��j������P�����Q�M��t�������賄���������@���_^[��  ;��r�����]���������������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������g��h�  ��$����w��P������Qy��j������Q�����R�M��Is������������������~���_^[��  ;�谆����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��*���   �H(�у�;��!����E�_^[���   ;�������]� ��������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������~��h�  ��$����u��P�������w��j������Q�����R�M���q�������葂������������_^[��  ;��P�����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M��Vk��h�  �������t��P�������8w��j �E�P������Q�M���k��������������������΁����������t�M�����M��K����E��M��;t��P�M�g����M��-����ER��P��p��XZ_^[��  ;��K�����]� �    ����   ,dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �BL�Ѓ�;�訃��_^[���   ;�蘃����]�������������������������U���  SVWQ�������E   ������Y�M��M��i��h�  ������Vs��P�������u��j �E�P������Q�M��Hj��������������������.�����������t�M�~����M�諍���E��M��r��P�M�Ǎ���M�荍���ER��P���cn��XZ_^[��  ;�諂����]� �   �����   �dat ����������������������������������������������������������������U���4  SVWQ�������M   ������Y�M��M��h��h�  �������&r��P�������ht��j �E�P������Q�M��i���������������������~����������t��ݝ ����M��{���݅ �����M��p}��ݝ����M��]���݅���R��P���0m��XZ_^[��4  ;��x�����]�   �����   �dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �B<�Ѓ�;��؀��_^[���   ;��Ȁ����]�������������������������U���,  SVWQ�������K   ������Y�M��M���f��h�  �������p��P��������r��j �E�P������Q�M��xg�������������������^}���������tǅ����    �M��ي����������M��e���������M�車�������R��P���k��XZ_^[��,  ;�������]Ë�   �����   �dat ����������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M��e��h�  ������Fo��P�������q��j �E�P������Q�M��8f��������������������|����������t�M�N����M�蛉���E�,�M������M���P�Q�P�Q�@�A�M��m����ER��P���Cj��XZ_^[��  ;��~����]� �   �����   �dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*���   �BP�Ѓ�;���}��_^[���   ;���}����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL���   �Ѓ�;��x}��_^[���   ;��h}����]�������������������������U����   SVWQ������9   ������Y�M���j�EP�M�Q�� ���R��*�HL���   �҃�;���|���M���P�Q�P�Q�@�A�E_^[���   ;���|����]� ����������������������������������������������U����   SVWQ������9   ������Y�M���j �EP�M�Q�� ���R��*�HL���   �҃�;��L|���M���P�Q�P�Q�@�A�E_^[���   ;�� |����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M��&b��h�  �������k��P�������n��j �E�P������Q�M��b��������������������x����������t�M�΀���M������E�,�M��t���M���P�Q�P�Q�@�A�M������ER��P�X!��f��XZ_^[��  ;��{����]� �   `!����   l!dat ����������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M���`��h�  ������j��P��������l��j �E�P������Q�M��xa��������������������^w����������t�M����M��ۄ���E�,�M��4~���M���P�Q�P�Q�@�A�M�譄���ER��P��"�e��XZ_^[��  ;���y����]� �   �"����   �"dat ����������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M��_��h�  ������Fi��P�������k��j �E�P������Q�M��8`��������������������v����������t�M�N~���M�蛃���E�,�M���|���M���P�Q�P�Q�@�A�M��m����ER��P��#�Cd��XZ_^[��  ;��x����]� �   �#����   �#dat ����������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M��f^��h�  �������h��P�������Hj��j �E�P������Q�M���^���������������������t����������tǅ���    �M��Y����������M�����������M��;��������R��P�%�c��XZ_^[��,  ;��Vw����]Ë�   %����    %dat ����������������������������������������������������������������������������U���  SVWQ�������B   ������Y�M����E�$�������x��h�  ��$����f��P�������h��j������P�����Q�M���b��������s���������)���_^[��  ;��[v����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�X�E�_^[��]� �������������������������������U���  SVWQ�������B   ������Y�M��EP�������_o��h�  ��$����e��P�������g��j������Q�����R�M���a��������r������������_^[��  ;��@u����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������l��h�  ��$�����d��P������!g��j������Q�����R�M��a���������q���������N��_^[��  ;��t����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q��*���   �H,�у�;���s���E�_^[���   ;���s����]� ��������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������j��h�  ��$����c��P�������e��j������Q�����R�M��_��������ap����������}��_^[��  ;�� s����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP��������i��h�  ��$����b��P������e��j������Q�����R�M���^��������o���������.}��_^[��  ;��`r����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������&i��h�  ��$�����a��P������Ad��j������Q�����R�M��9^���������n���������n|��_^[��  ;��q����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP��������j��h�  ��$����?a��P������c��j������Q�����R�M��y]��������!n���������{��_^[��  ;���p����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M���V��h�  ������`��P��������b��j �E�P������Q�M��xW��������������������^m����������t�M�u���M���z���E�,�M��4t���M���P�Q�P�Q�@�A�M��z���ER��P��,�[��XZ_^[��  ;���o����]� �   �,����   �,dat ����������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M��U��h�  �������F_��P�������a��j �E�P������Q�M��8V��������������������l����������tǅ���    �M��y���������M��%~��������M��{y�������R��P��-�NZ��XZ_^[��,  ;��n����]Ë�   �-����   �-dat ����������������������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M��fT��h�  �������^��P�������H`��j �E�P������Q�M���T���������������������j����������tǅ���    �M��Yx���������M���|��������M��;x�������R��P�/�Y��XZ_^[��,  ;��Vm����]Ë�   /����    /dat ����������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M���x���E�}�t�}�t�}�tǅ$���    �
ǅ$���   ��$���_^[���   ;��l����]���������������������������������U���  SVWQ�������B   ������Y�M��EP�������Vc��h�  ��$����/\��P������q^��j������Q�����R�M��iX��������i���������v��_^[��  ;���k����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������/e��h�  ��$����o[��P������]��j������Q�����R�M��W��������Qh����������u��_^[��  ;��k����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������od��h�  ��$����Z��P�������\��j������Q�����R�M���V��������g���������u��_^[��  ;��Pj����]� ����������������������������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;���i��_^[���   ;���i����]������������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;��mi��_^[���   ;��]i����]������������������������������U����   SVW��@����0   �����󫡘*�H�􋑘   ��;��i��_^[���   ;���h����]����������������������U����   SVW��@����0   �����󫡘*�H�􋑜   ��;��h��_^[���   ;��h����]����������������������U����   SVW��@����0   �������E�Q��*�B���   �у�;��;h���E�     _^[���   ;��"h����]�����������������������������������U����   SVW��@����0   �������EP��*�Q���   �Ѓ�;��g��_^[���   ;��g����]������������������������������U����   SVW��4����3   �������ja���E��}� u3��_��EP�MQ�UR�E�P��*�Q���  �Ѓ�;��/g����u+�}� t��E�P��*�Q@�B�Ѓ�;��g���E�    �E�_^[���   ;���f����]����������������������������������������������U����   SVW��@����0   �������EPj �MQ�a����P�UR�EP��*�Q���  �Ѓ�;��ff��_^[���   ;��Vf����]���������������������������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q���   �Ѓ�;��e��_^[���   ;��e����]����������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP��*�Q���   �Ѓ�;��e��_^[���   ;��e����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�BL�Ѓ�;��d��_^[���   ;��d����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�BP�Ѓ�;��+d��_^[���   ;��d����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�HL�QT�҃�;��c��_^[���   ;��c����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL��  �у�;��4c��_^[���   ;��$c����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL���   �у�;��b��_^[���   ;��b����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�BX�Ѓ�;��;b��_^[���   ;��+b����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�QL�B\�Ѓ�;��a��_^[���   ;��a����]� �����������������������������U���T  SVWQ�������U   ������Y�M��e[���E�}� u3��  �E�    �E�    �E�    �M��G���M��v���E�E��E��E��EPh]  �M��JV��j j �E�P�M���t����u��   �M��HF���E���E��Eȃ}� ��   �M���q���E��EȉE��E�Ph�   ��K������u�   �}� u�~j �M��.E���Eԃ}� u�i�E�P�M��N���E�P�!d�����}� t��E�P��*�Q@�B�Ѓ�;��X`���E�    �`����E쉅�����M��Df���M��'I���������W�}� t��E�P��*�Q@�B�Ѓ�;��`���E�    �E�P�c����ǅ����    �M���e���M���H��������R��P��<�kK��XZ_^[��T  ;��_����]� �   �<����   �<����   �<cd ctr �����������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*���   �M��B��;��!^��_^[���   ;��^����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M����   ��;��]��_^[���   ;��]����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M��B<��;��(]��_^[���   ;��]����]� ����������������������U����   SVWQ��4����3   ������Y�M���*���   ��M��B(��;��\��_^[���   ;��\����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�B`�Ѓ�;��K\��_^[���   ;��;\����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�Bd�Ѓ�;���[��_^[���   ;���[����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL�Hh�у�;��g[��_^[���   ;��W[����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL��D  �Ѓ�;���Z��_^[���   ;���Z����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL�Bl�Ѓ�;��{Z��_^[���   ;��kZ����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BL���   �у�;��Z��_^[���   ;���Y����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M$�H��h�Dh Dh�Ch`C�E��HQ�U R�EP�MQ���E�$�UR�E��HQ�U�R��*�HL���   �҃�4;��<Y��_^[���   ;��,Y����]�  ������������������������������������������U����   SVW��@����0   ������E���M���;���X��_^[���   ;��X����]��������������������������U����   SVW��@����0   �������EP�M��M�B��;��dX��_^[���   ;��TX����]���������������������U����   SVW��@����0   �������EP�MQ�U��M�P��;�� X��_^[���   ;���W����]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�M��M�B��;��W��_^[���   ;��xW����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QL���   �Ѓ�;��W��_^[���   ;��W����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�QL��   �Ѓ�;��V��_^[���   ;��V����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ��*�BL�M���H  ��;��V��_^[���   ;��V����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���*�PL��M���L  ��;��U��_^[���   ;��U����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�QL�M���P  ��;��(U��_^[���   ;��U����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�QL�M���T  ��;��T��_^[���   ;��T����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�HL���   �҃�;��5T��_^[���   ;��%T����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�QL���   �Ѓ�;��S��_^[���   ;��S����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�BL��   �у�;��(S��_^[���   ;��S����]� ��������������������������������������U���  SVW�������B   ������M��g���M���X���} t�M���f����u"ǅ����   �M��\6���M��X���������Qj�M��f��P�M��L���M��f���E�E�E��E�Ph=���c=����������M��	6���M��HX�������R��P�HJ��=��XZ_^[��  ;��R����]�   PJ����   oJ����   hJactive mu ������������������������������������������������������������������������������U���  SVW�������B   ������M��Hf���M��W���} t�M��e����u"ǅ����   �M��5���M��KW���������Qj�M��]e��P�M�K���M��Le���E�E�E��E�Ph<���<����������M��4���M���V�������R��P��K�<��XZ_^[��  ;���P����]�   �K����   �K����   �Kactive mu ������������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR��*�HL���   �҃�;��P��_^[���   ;���O����]�����������������������U����   SVW��@����0   �������EP�MQ��*�BL���   �у�;��O��_^[���   ;��O����]��������������������������U����   SVW��@����0   �������EP�MQ��*�BL���   �у�;��)O��_^[���   ;��O����]��������������������������U����   SVW��@����0   �����󫡘*�HL��  ��;���N��_^[���   ;��N����]����������������������U����   SVW��@����0   �����󫡘*�HL��@  ��;��eN��_^[���   ;��UN����]����������������������U����   SVWQ��(����6   ������Y�M�j\�f   ���E�}� t	�E�x\ u���EP�M�Q�U�B\�Ѓ�;���M��_^[���   ;���M����]� �����������������������������U����   SVW��@����0   ������h�/�EPh^� �_����_^[���   ;��hM����]�������������������������U����   SVWQ��4����3   ������Y�M��\8���M���E�_^[���   ;��M����]�����������������������������U����   SVW��@����0   �����󫡘*���   �􋑈   ��;��L��_^[���   ;��L����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�P��O�����E��     _^[���   ;��4L����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@���E�@8���E�@<~��E�@@��E�@D��E�@H���E�@L���E�@P*��E�@l��E�@X���E�@\���E�@`��E�@dɘ�E�@TĘ�E�@h���E�@p���E�@tΘ�E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������������U���h  SVW�������Z   ������j h�   ��\���P�`K����j �EP�MQ�UR�EP��\���Q�]P�����E �E�h�   ��\���P�MQ�URj�O?����R��P�pV�1��XZ_^[��h  ;���E����]Ë�   xV\����   �Vnp ���������������������������������������������������������U����   SVW��@����0   ������EP�M���   Q�UR�[����_^[���   ;��TE����]���������������������U���  SVWQ��\����i   ������Y�M���.���M���E��8 u��   �EP��l�����Y��j h����������N��P��������Y��j j���l���Q������R������P�Z����P������Q�=����P�����R�=����P�E����*��������؈�c����������1���������1���������1���������1����������W����l����1����c�����t�E�P��,�����E�_^[�Ĥ  ;��D����]� ��������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�p:�����M���E�_^[���   ;��eC����]� �������������������U����   SVWQ��4����3   ������Y�M��E�P��+����_^[���   ;��C����]�����������������������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��M�BG���E_^[���   ;��@����]� ����������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����  SVW��(����v   ������ǅ ���    �}( uǅ0���    �M�JS����0����!  �E�    �M�zJ������  �M��?���M���1������   �EP��H����}T���� ���j h���������yI���� ���P��l����QT���� ���j j���H���Q��l���R������P�U������ ���P������Q�'8������ ���P������R�8������ ��� P�M���%�����J%����uǅ(���   �
ǅ(���    ��(�����?����� ����� t�� ���ߍ�������+���� �����t�� ���������+���� �����t�� ������������+���� �����t�� ������l����+���� �����t�� �����������Q���� �����t�� ������H����n+����?�����t(�E(P�M$Q�M��+0��P�UR�EP�MQ�gP�����E��M��#J���!�E(P�M$Qj �UR�EP�MQ�<P�����E��E�������M�$Q�������R��P��^�7)��XZ_^[���  ;��=����]ÍI    �^����   �^icon �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��'K�������_^[���   ;��k<����]����������������������������U���  SVW��x����b   ������} u3��   j h�   ��<���P�A�����E��\����E��|����E�E��E��<���ǅ@������E�%��E���E����E����E�,��E����E�ԡh�   ��<���P�MQ�URj��4����R��P��`�('��XZ_^[�Ĉ  ;��p;����]�   �`<����   anp �������������������������������������������������������������������������U���  SVW��x����b   ������j h�   ��<���P��?����ǅ\���    �E��|���h�   ��<���P�MQ�URj��3����R��P��a�>&��XZ_^[�Ĉ  ;��:����]Ë�   �a<����   �anp ��������������������������������������������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`�����������U����   SVW��@����0   �����󫡘*�H���   ��;��9��_^[���   ;��9����]����������������������U����   SVW��@����0   �������E�Q��*�B���   �у�;��+9���E�     _^[���   ;��9����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q���   �Ѓ�;��8��_^[���   ;��8����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B���   �у�;��48��_^[���   ;��$8����]� ����������������������������������U����   SVW��@����0   �����󫡘*�H����;���7��_^[���   ;��7����]��������������������������U����   SVW��@����0   �������E�Q��*�B�H�у�;��^7���E�     _^[���   ;��E7����]��������������������������������������U����   SVW��@����0   �������E�Q��*�B�H�у�;���6���E�     _^[���   ;���6����]��������������������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q��*�B���   �у�;��L6�����E��������� �����@�������_^[���   ;��6����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;��5��_^[���   ;��5����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�H\�у�;��75��_^[���   ;��'5����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�H���   �҃�;��4��_^[���   ;��4����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B�HX�у�;��4��_^[���   ;��4����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B �Ѓ�;��3��_^[���   ;��3����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B���   �у�;��(3��_^[���   ;��3����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q�B�Ѓ�;��2��_^[���   ;��2����]� �����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ��*�B��   �у�;��2��_^[���   ;��2����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q�M��B$��;��1��_^[���   ;��1����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B�H(�у�;��1��_^[���   ;��1����]� �������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P��*�Q�B`�Ѓ�(;��0��_^[���   ;��w0����]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B�H,�у�;���/��_^[���   ;���/����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��<����P�M���?����Pj j �E�P��*�Q�B4�Ѓ� ;��c/��_^[���   ;��S/����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q��*�B�H4�у� ;���.��_^[���   ;��.����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H�Q@�҃�;��T.��_^[���   ;��D.����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�HD�у�;���-��_^[���   ;���-����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�BL�Ѓ�;��[-��_^[���   ;��K-����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�BL�Ѓ�;���,��_^[���   ;���,����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�BP�Ѓ�;��{,��_^[���   ;��k,����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�HT�у�;��,��_^[���   ;���+����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�HT�у�;��+��_^[���   ;��w+����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���   �҃�;��+��_^[���   ;���*����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P��*�Q���   �Ѓ�;��y*��P�M��*���� ����#5���E_^[���   ;��R*����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�Bh�Ѓ�;���)��_^[���   ;���)����]����������������������������U����   SVW��0����4   ������h��D��Ph�/h�   �(2������8�����8��� t��8����7����0����
ǅ0���    ��0���_^[���   ;��<)����]���������������������������������������������U����   SVW��$����7   ������E�8 t?�E���8�����8�����,�����,��� tj��,����5����$����
ǅ$���    �E�     _^[���   ;��(����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����E��t�E�P������E�_^[���   ;��
(����]� ������������������������U����   SVWQ��4����3   ������Y�M��M����� ���M���,���E�_^[���   ;��'����]��������������������U����   SVWQ��(����6   ������Y�M��M���/���E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��&'����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M��$���M������_^[���   ;��&����]�����������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��a&����]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E����Xp�E��@x�����E��@|   _^[��]������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	�-���E��     �E��x` t�E���`P�����_^[���   ;��I%����]������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 th��H��P������E��x` th��H��P�r�����M�����M���)���E�P�M���dQ�U��BxP�MQ�U���`R�.�����M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�������E��@|�   �E��xd ��   �E���pP�M���hQ�UR��!������u(�E��@h    �E����Xph��H��P������EP�M�����.��j j j�E���P�M��	�M+���U��B|�E��x|t�M������E��@|��E��@x�����E��@|_^[���   ;��z#����]� ������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��$���M���'��_^[���   ;��"����]��������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	��)���U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;���!����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap��E��xd t�E��@h��E��x|u�   �3�_^[��]� ��������������������������������U����   SVW��@����0   �����󫡘*�H����;��� ��_^[���   ;��� ����]��������������������������U����   SVW��@����0   �������E�Q��*�B�H�у�;��~ ���E�     _^[���   ;��e ����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q��*�B�H�у� ;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B�H�у�;��g��_^[���   ;��W����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H�Q�҃�;��t��_^[���   ;��d����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��r�����M��h���H �G@��;�����_^[���   ;�������]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��������M������H �GD��;��Z��_^[���   ;��J����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M��`���xH u3��#�M��N�����M��D�����H �FH��;�����_^[���   ;������]�������������������������������������U����   SVWQ��4����3   ������Y�M��M������xL u3��/��EP�MQ�UR�M�������M�����H �GL��;��(��_^[���   ;������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M��0���xP u����3��EP�MQ�UR�EP�M�������M�����H �WP��;����_^[���   ;��s����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M�����xT u����+��EP�MQ�M��s�����M��i���H �WT��;�����_^[���   ;�������]� �����������������������������������������U���  SVWQ�������C   ������Y�M��} t<�M��� ����E�P�M��� �����M��� ���H �WL��;��T���M��M��;���} t?������� ��P�M��/���������-���M�� ���@@�EЃ}� t�E�P�M�/��R��P������XZ_^[��  ;�������]� �I    ������   ��bc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������x` u� }  �'��EP�M��������M������H �W`��;����_^[���   ;������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��������M������H �WH��;����_^[���   ;������]� ��������������������������������U����   SVWQ��(����6   ������Y�M�j�EP�$���������P�M��*-���E�M�V(��;E��M�u$��;E�~������3��EP�MQ�UR�EP�M��M������M��C����H �WD��;�����_^[���   ;������]� ���������������������������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M������xP u������;��EP�MQ�UR�EP�MQ�UR�M��Q������M��G����H �GP��;�����_^[���   ;������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�������xT u������+��EP�MQ�M��������M������H �WT��;��)��_^[���   ;������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��0����xX u�'��EP�M��������M������H �WX��;����_^[���   ;������]� ��������������������������������U����   SVW�� ����8   ������M�����E�P�MQ��#������t�}� u3���E�P�M�Q�U�R�E�P�M�����R��P���� ��XZ_^[���   ;�������]ÍI    ������   ��dat ����������������������������������������������������U����   SVWQ������<   ������Y�M��M�����M�������uh��L��P�������3��   �E�    ��E�P�M�Q�UR�E�P��*�Q���   �Ѓ�;������u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�'���͍E�P�
�����   R��P�Ԉ�F���XZ_^[���   ;������]�    ܈����   ������   �arr count ����������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M�8����M��h����uh��P��P�u�����3��   �E�    ��E�P�M�Q�UR�E�P��*�Q���   �Ѓ�;������u3��i�}� u3��_�E�    �	�Eԃ��EԋE�;E�}4�EԋM��<� t�EԋM���������u�ϋEԋM���R�M�;��뻍E�P�������   R��P�p�����XZ_^[���   ;�������]�    x�����   ������   ��arr count ��������������������������������������������������������������������������������������U����   SVW��@����0   �����󫡘*�H��   ��;��5��_^[���   ;��%����]����������������������U����   SVW��@����0   �������E�Q��*�B��$  �у�;������E�     _^[���   ;������]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��*�B��(  �у�;��D���E�_^[���   ;��1����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��*�B��,  �у�;�����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ��*�B��,  �у�;��D�������_^[���   ;��-����]� ���������������������������U����   SVW��@����0   �����󫡘*�H��0  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡘*�H��4  ��;��u��_^[���   ;��e����]����������������������U����   SVWQ��0����4   ������Y�M��} t�M�/	����0����
ǅ0���    ��0���P�M�Q��*�B��8  �у�;�����_^[���   ;�������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B��<  �у�;��T��_^[���   ;��D����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q��@  �Ѓ�;�����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H��D  �҃�;��Q��_^[���   ;��A����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B��H  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R��*�H��L  �҃�;��N��P�M������ �������E_^[���   ;��'����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q��T  �Ѓ�;��
��_^[���   ;��
����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q��P  �Ѓ�;��H
��_^[���   ;��8
����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B��X  �у�;���	��_^[���   ;���	����]� ����������������������������������U����   SVW��@����0   �����󫡘*�H��\  ��;��e	��_^[���   ;��U	����]����������������������U����   SVW��@����0   �������E�Q��*�B��`  �у�;������E�     _^[���   ;�������]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�H��d  �҃�;��e��_^[���   ;��U����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R��*�H��h  �҃�;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��G���_^[���   ;��]����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;������]������������������U����   SVWQ��4����3   ������Y�M��EP�M�����_^[���   ;������]� ���������������������������U����   SVWQ��4����3   ������Y�M��M��c���_^[���   ;��Q����]������������������U����   SVWQ��4����3   ������Y�M��E�� �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��*����E��t�E�P�������E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]��������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;�����������
ǅ���    �E�    _^[���   ;������]������������������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M���  ��;��=��_^[���   ;��-����]������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M���(  ��;�����_^[���   ;������]������������������������������U����   SVWQ������<   ������Y�M������P��*�Q�M���   ��;��U��P�M�<������������E_^[���   ;��.����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���*�P��M���$  ��;����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP�MQ��*�B��  �у�;��I��_^[���   ;��9����]��������������������������U����   SVW��@����0   �������EP��*�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �����󫡘*�H��  ��;��u��_^[���   ;��e����]����������������������U����   SVW��@����0   �������EP�MQ�UR��*�H���  �҃�;����_^[���   ;��� ����]�����������������������U����   SVW��@����0   �������EP�MQ��*�B��x  �у�;�� ��_^[���   ;�� ����]��������������������������U����   SVW��@����0   �������EP��*�Q��|  �Ѓ�;��- ��_^[���   ;�� ����]������������������������������U����   SVWQ��0����4   ������Y�M��E�M��;t3���   �E�x uN�E�8 uF�E�x u=�E��x u�M��9 u�U��z uǅ0���   �
ǅ0���    ��0����   �R�E��x uI�E��8 uA�E��x u8�E�x u�M�9 u�U�z uǅ0���   �
ǅ0���    ��0����M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� �������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M����������_^[���   ;��&�����]� ��������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M��b����8 t��E�_^[���   ;�������]����������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M�������8 t(�E�P�M�����P�M�Q�M��������������t�뾃} t�E�M��}� ~�E�P�M������8 uǅ$���   �
ǅ$���    ��$���_^[���   ;��������]� �����������������������������������������������������������U����   SVW��4����3   ������j�k   ���E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;��.���_^[���   ;�������]�������������������������������U����   SVW��@����0   ������h\/�EPhD �	����_^[���   ;�������]�������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u���E�P�M�Q\�҃�;��C����E�_^[���   ;��0�����]���������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;������EP�M��[
���E�_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;������EP�M��,����E�_^[���   ;��������]� ����������������������������������U����   SVWQ������;   ������Y�M�j\�������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;��s����EP������y���P�M������E�_^[���   ;��H�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;�������EP�M�������EP�M�������E�_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;������EP�M��,����EP�M��$����EP�M������E�_^[���   ;��������]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�������E�}� t	�E�x` u���E�P�M�Q`�҃�;��S���_^[���   ;��C�����]������������������������������������U����   SVWQ��(����6   ������Y�M�jd��������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jh�f������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;��/���_^[���   ;�������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jl��������E�}� t	�E�xl u���E�P�M�Ql�҃�;�����_^[���   ;�������]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��d���_^[���   ;��T�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u�`/���EP�M�Q�U�Bp�Ѓ�;������_^[���   ;�������]� ����������������������������������������U����   SVWQ������:   ������Y�M�jt�f������E�}� t	�E�xt uh`/�M�����E�:��EP�M�Q�����R�E�Ht�у�;�����P�M����������*����E_^[���   ;��������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�������E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;��\����E�_^[���   ;��I�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jx��������E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�V������E�}� t	�E�x| u�   �#��E�P�MQ�U�B|�Ѓ�;����������_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��4����3   ������j�{������E��}� t	�E��x u3���E���H��;��M���_^[���   ;��=�����]������������������������������U����   SVW��4����3   ������E�8 u�?j��������E��}� t	�E��x u�!��EP�M��Q�҃�;������E�     _^[���   ;�������]��������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j�L������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;�����_^[���   ;��������]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��m���_^[���   ;��]�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;������_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �f������E�}� t	�E�x  u3����E�P�M�Q �҃�;��1���_^[���   ;��!�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;�����_^[���   ;�������]����������������������������������U����   SVWQ��(����6   ������Y�M�j(�F������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;�����_^[���   ;��������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;��i���_^[���   ;��Y�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;������_^[���   ;�������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j4�f������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��1���_^[���   ;��!�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8��������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;�����_^[���   ;�������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�&������E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;������_^[���   ;��������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jD�������E�}� t	�E�xD u3����E�P�M�QD�҃�;��a���_^[���   ;��Q�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� u���EP�M�Q�U�BH�Ѓ�;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jL�v������E�}� u3����EP�M�Q�U�BL�Ѓ�;��F���_^[���   ;��6�����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�jP��������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;�����_^[���   ;�������]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�V������E�}� u3����E�P�M�QT�҃�;��*���_^[���   ;�������]���������������������������U����   SVWQ��(����6   ������Y�M�jX��������E�}� u���EP�M�Q�U�BX�Ѓ�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;�� ���_^[���   ;��������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��X���_^[���   ;��H�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;������_^[���   ;�������]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��0���_^[���   ;�� �����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;�������]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��
���_^[���   ;��������]� ����������������������������������������U����   SVW������9   ������h�   �������E��}� u�M�����E�9��EP�� ���Q�U����   �Ѓ�;��i���P�M������� ���������E_^[���   ;��B�����]���������������������������������������������������U����   SVWQ������?   ������Y�M�h�   ��������E�}� t�E샸�    uj ����������P�M�����E�9��EP�����Q�U�M����   ��;�����P�M��������������E_^[���   ;��c�����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;������_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3����EP�U�M����   ��;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;��x���_^[���   ;��h�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����E�M����   ��;��<���_^[���   ;��,�����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;�����_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u���EP�U�M����   ��;������_^[���   ;��������]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��@���_^[���   ;��0�����]� ����������������������������������������������U����   SVWQ������9   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�M����   ��;������E��E�_^[���   ;�������]���������������������������������������U����   SVWQ��(����6   ������Y�M���E�P��*���   �BX�Ѓ�;������E�}� u3���EP�MQ�M��g���_^[���   ;��������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H|�Q�҃�;��t���_^[���   ;��d�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P��*���   �BX�Ѓ�;�������E�}� u3���EP�MQ�M��K���_^[���   ;��������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H|�Q8�҃�;��T���_^[���   ;��D�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q��*�B�H�у�;�������U��B�E�_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q��*�B�H�у�;��C����U��B_^[���   ;��-�����]������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��E��HQ�UR�EP�M��R��*�H�Q�҃�;������M��A�   _^[���   ;�������]� ���������������������������������U����   SVW��<����1   ������E��<�����<���t��E�x/�E�t/�   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$�,��   �]  �|/���|/�=|/��   �EP������=�.  }
������&  �} u
������  h�T��Ph�/j��������� ����� ��� t�� �������������
ǅ���    ������p/�=p/ t�EP�p/������   �   �EP�MQ��������u����   �   �|������u�|/���|/u\�����A����=p/ t?�p/��8�����8�����,�����,��� tj��,����R���������
ǅ���    �p/    �   ����_^[���   ;��5�����]Ð���������x�����������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M����]����z	���]�x�]����Au	�x�]�E�h�h���$��������E���E��h�X�M������E�_^[���   ;��������]� ��������������������������������������������U����   SVWQ�� ����8   ������Y�M����]����Azǅ$���   �
ǅ$���    ���]����Azǅ ���   �
ǅ ���    ��$���3�;� ������M���E�$�.������h���$�ӿ�����E�����E�$�������h���$詿�����E��X�E����X����Auh��X��P荺�����E����X�}� u�E�� ���M���M��5����E�_^[���   ;�������]� ��������������������������������������������������������������������������������U����   SVW��@����0   ��������E�$�g�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X�E����X����Auh��\��P�Q������E����X_^[���   ;�������]� ���������������������������������U����   SVWQ��,����5   ������Y�M����]����Auh��`��P�͸�������]�E�� �M���$製�����M����A�$ݝ,���艽����ܽ,������$�u������U�����E�$�_������E��X�M��*���_^[���   ;�������]� ��������������������������������������������������������U���0  SVWQ�������L   ������Y�M��E���� �$�������]�E����@�$��������]���]�����At��]�����Au�E�����E����X�U  � �]�����Auz� �]�����Auj�E�������E��E�������E��}� u�E�����E����X�8�E���}��U��E��E��E��E��}� u��E��E��8�M���E��E��x�M��Y��   ���E��$���E��$�������=��]����]�����Au.�E��M��]��E��M��]؋E�� �M��M���E��@�M��M��Y���]�����Au���]؋E����X���E��$���E��$��������]��E��]��E��]��h�]�����A{ǋE�� �u�M���E��@�u�M��Y_^[��0  ;��s�����]������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������E�]����Au�E��E_^[��]�����������������������U����   SVW��@����0   ������E���M�B��;��h���_^[���   ;��X�����]�������������������������U����   SVW��@����0   ������E���M�B��;�����_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M��E��  �E��@    ��h`��E�Ph��h���*�QP��Ѓ�;��z����M��A�E�_^[���   ;��a�����]����������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVW��@����0   ������E���M�B��;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M��M��N����E��t�E�P�L������E�_^[���   ;��J�����]� ������������������������U����   SVWQ��4����3   ������Y�M��E��  �E��x u!��E��HQ��*�BP�H�у�;������_^[���   ;��������]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��+��j �EP�MQ�U��BP��*�QP�B�Ѓ�;��A���_^[���   ;��1�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��x t$��EP�M��QR��*�HP�Q�҃�;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M��E��x t$��EP�M��QR��*�HP�Q�҃�;��<���_^[���   ;��,�����]� ��������������������������U����   SVW��@����0   �����󫡘*�HP�􋑈   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������EP��*�QP���   �Ѓ�;��m���_^[���   ;��]�����]������������������������������U����   SVW��@����0   �����󫡘*�HP��QP��;�����_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP��*�QP�BT�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��8 u�I��E��Q��*�BP�HL�у�;��������E��Q��*�BP�H<�у�;������E��     _^[���   ;�������]���������������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M����P�M��+���_^[���   ;�� �����]� ������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��(����6   ������Y�M��E��8 t3��E��Q��*�BP�H<�у�;��q����E��     �E��@    �E��M�H��h`��EPh��h��MQ�UR��*�HP�Q8�҃�;��!����M���E�    �	�E���E�E�;E}z�E�M���z u7�E�M���B   �E�M����BP��*�QP�B�Ѓ�;�������E�P�M��R��*�HP�Q@�҃�;������M�U���A�u����E�3Ƀ8 ����_^[���   ;��k�����]� �����������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H}��E�P�M��R��*�HP�Q@�҃�;������E�}� t*��j �EPj�M�Q��*�BP�H�у�;��s�����u$��E��Q��*�BP�HL�у�;��O���3��
�m����   _^[���   ;��1�����]� ���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E��Q��*�BP�HD�у�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���E��Q��*�BP�HH�у�;��9���_^[���   ;��)�����]��������������������������U����   SVWQ��4����3   ������Y�M���E��Q��*�BP�HL�у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ������_^[���   ;��K�����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�������E��}� u3��5�M��ʮ���E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;��Y�����]������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E��     �E��@    �E��@   �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��} u�4�} t�EP�M����� �} t�EP�M�|�����E�P�M�n���_^[���   ;��M�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M��B@��;��ؽ��_^[���   ;��Ƚ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M��BD��;��h���_^[���   ;��X�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M��Bd��;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M��Bh��;�苼��_^[���   ;��{�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B@�M��Pl��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B@�M��Pp��;�藻��_^[���   ;�臻����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP��*���   �M����   ��;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*���   �M����   ��;�葺��_^[���   ;�聺����]� �������������������������������U����   SVWQ��4����3   ������Y�M���*�P@��M��Bt��;�� ���_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���*�P@��M��Bx��;�谹��_^[���   ;�蠹����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M��B|��;��;���_^[���   ;��+�����]� �������������������������U����   SVWQ��4����3   ������Y�M���*�P@��M����   ��;��͸��_^[���   ;�轸����]������������������������������U����   SVWQ��4����3   ������Y�M���*���   ��M��Bt��;��]���_^[���   ;��M�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M����   ��;�����_^[���   ;��ط����]� ����������������������U����   SVWQ��4����3   ������Y�M���*�P@��M����   ��;��}���_^[���   ;��m�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M����   ��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*�Q@�M����   ��;�茶��_^[���   ;��|�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P@�M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*�P@�M����   ��;�葵��_^[���   ;�聵����]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P��*�Q@�B�Ѓ�;������E�E�#Et�E��#E�E��	�E�E�E��E�P�M�Q��*�B@�H�у�;��ش��_^[���   ;��ȴ����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QH���   �Ѓ�;��X���_^[���   ;��H�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B@�HL�у�;�����_^[���   ;��׳����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q@�BH�Ѓ�;��k���_^[���   ;��[�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q@�B�Ѓ�;�����_^[���   ;��߲����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B@�H�у�;��w���_^[���   ;��g�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H@�Q�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�B@�H �у�;��w���_^[���   ;��g�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*���   �M��P��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*���   �M��B��;��q���_^[���   ;��a�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*���   �M��B ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP��*���   �M����   ��;��i���_^[���   ;��Y�����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR��*���   �M���D  ��;��ޮ��_^[���   ;��ή����]� ����������������������������U����   SVWQ��4����3   ������Y�M���E P���E�$�MQ�UR�EP�MQ��*���   �M����   ��;��L���_^[���   ;��<�����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ��*���   �M����   ��;�赭��_^[���   ;�襭����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���*���   ��M��B$��;��=���_^[���   ;��-�����]������������������������������U����   SVW��@����0   �����󫡘*�H@��Q0��;��ج��_^[���   ;��Ȭ����]�������������������������U����   SVW��@����0   �������j�EPj ��*�Q@�B4�Ѓ�;��l���_^[���   ;��\�����]�����������������������������U����   SVW��@����0   �������j�EPh   @��*�Q@�B4�Ѓ�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQj ��*�B@�H4�у�;�芫��_^[���   ;��z�����]���������������������������U����   SVW��@����0   �����󫡘*�H|����;��)���_^[���   ;�������]��������������������������U����   SVW��@����0   ������E�8 t ��E�Q��*�B|�H�у�;�趪���E�     _^[���   ;�蝪����]������������������������������U����   SVW��@����0   �����󫡘*�H|��Q ��;��H���_^[���   ;��8�����]�������������������������U����   SVW��@����0   ������E�8 t ��E�Q��*�B|�H(�у�;��֩���E�     _^[���   ;�轩����]������������������������������U����   SVW��@����0   �����󫡘*�H@��Q0��;��h���_^[���   ;��X�����]�������������������������U����   SVW��@����0   ������E�8 t ��E�Q��*�B@�H�у�;�������E�     _^[���   ;��ݨ����]������������������������������U����   SVW��@����0   �������EP��*�Q@���   �Ѓ�;��}���_^[���   ;��m�����]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q��*�B@�H�у�;������E�     _^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�QH���   �Ѓ�;�舧��_^[���   ;��x�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BH��d  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q �BH�Ѓ�;�蔦��_^[���   ;�脦����]�������������������������������������U����   SVW��4����3   ������}qF t�1�E�E��}� u�#�EP�M��*����E�P�MQ�M�x������ݶ��_^[���   ;�������]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B�M��Pp��;�臥��_^[���   ;��w�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q@�B,�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���*�P@��M��BT��;�蠤��_^[���   ;�萤����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q@�M��BX��;��+���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ��*�B@�M��P\��;�跣��_^[���   ;�解����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���*�P@��M��B`��;��@���_^[���   ;��0�����]���������������������������������U����   SVW��@����0   �������EP�MQ��*�B��T  �у�;��ɢ��_^[���   ;�蹢����]��������������������������U����   SVW��@����0   ������h��hE  �M�ۍ����������Ph��hE  �M迍��������P��*�H��T  �҃�;��.���_^[���   ;�������]�����������������������������������������������U����   SVWQ��(����6   ������Y�M�j�v   ���E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;�艡��_^[���   ;��y�����]� ���������������������������������������U����   SVW��@����0   ������h�/�EPh^� �Y�����_^[���   ;�������]�������������������������U����   SVWQ��(����6   ������Y�M�j�v������E�}� t	�E�x u3����E�P�M�Q�҃�;�葠��_^[���   ;�聠����]����������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u���� ��EP�MQ�U�R�E�H�у�;������_^[���   ;�������]� ��������������������������������������U���h  SVWQ��������   ������Y�M�j�F������E�}� t	�E�x u�M�m����E�2��EP�M�Q������R�E�H�у�;��M����b   ���}�E_^[��h  ;��.�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M������M���`�����M����   �ע���M���   �ɢ���E���ݘ�  �E�_^[���   ;�茞����]���������������������������������������������U���L  SVWQ�������S   ������Y�M��M��o����M����d����M���0�Y����M���H�N��������$�����$�����$�����������M����P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������А���M������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������腐���M���0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������:����M���H���P�Q�P�Q�P�Q�P�Q�@�A�E�_^[��L  ;��Ԝ����]�����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��E��E��E�X�E��E�X�E�_^[��]� �����������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u� ��EP�MQ�U�R�E�H�у�;�諛��_^[���   ;�蛛����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u�$��EP�MQ�UR�E�P�M�Q�҃�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��(����6   ������Y�M�j �V������E�}� t	�E�x  u3��$��EP�MQ�UR�E�P�M�Q �҃�;��e���_^[���   ;��U�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u3����EP�M�Q�U�B$�Ѓ�;��͙��_^[���   ;�轙����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x( u�(��EP�MQ�UR�EP�M�Q�U�B(�Ѓ�;��#���_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j,�v������E�}� t	�E�x, u��� ��EP�MQ�U�R�E�H,�у�;�艘��_^[���   ;��y�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j0��������E�}� t	�E�x0 u3��)����E�$�EP�MQ�U�R�E�H0�у�;������_^[���   ;��З����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4�&������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��A���_^[���   ;��1�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u���E�P�M�Q8�҃�;�賖��_^[���   ;�裖����]������������������������������������U���@  SVWQ�������P   ������Y�M�jD�������E�}� t	�E�xD u�M�T����E�.��E�P������Q�U�BD�Ѓ�;������   ���}�E_^[��@  ;�������]� ������������������������������������������������U����   SVWQ��(����6   ������Y�M�jH�F������E�}� t	�E�xH u���EP�M�Q�U�BH�Ѓ�;��_���_^[���   ;��O�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jL�������E�}� t	�E�xL u������EP�M�Q�U�BL�Ѓ�;��̔��_^[���   ;�輔����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�jP�������E�}� t	�E�xP u���EP�M�Q�U�BP�Ѓ�;��/���_^[���   ;�������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jT�������E�}� t	�E�xT u���EP�M�Q�U�BT�Ѓ�;�蟓��_^[���   ;�菓����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jX��������E�}� t	�E�xX u3��4��E P�MQ�UR�EP�MQ�UR�EP�M�Q�U�BX�Ѓ� ;������_^[���   ;�������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j`�F������E�}� t	�E�x` u3����E�P�M�Q`�҃�;��a���_^[���   ;��Q�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jd�������E�}� t	�E�xd u3����EP�M�Q�U�Bd�Ѓ�;��͑��_^[���   ;�轑����]� �������������������������������������������U����   SVWQ������:   ������Y�M�jh�������E�}� t	�E�xh u�M�0����E�:��EP�M�Q�����R�E�Hh�у�;�����P�M�|��������/����E_^[���   ;��������]� ����������������������������������������������������U����   SVWQ��(����6   ������Y�M�jp�F������E�}� t	�E�xp u������E�P�M�Qp�҃�;��`���_^[���   ;��P�����]���������������������������������U����   SVWQ��(����6   ������Y�M�jl�������E�}� t	�E�xl u������E�P�M�Ql�҃�;��Џ��_^[���   ;��������]���������������������������������U����   SVWQ��(����6   ������Y�M�jt�&������E�}� t	�E�xt u3����E�P�M�Qt�҃�;��A���_^[���   ;��1�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jx�������E�}� t	�E�xx u���EP�M�Q�U�Bx�Ѓ�;�诎��_^[���   ;�蟎����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j|�������E�}� t	�E�x| u���E�P�M�Q|�҃�;��#���_^[���   ;�������]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u���E�P�M싑�   �҃�;�芍��_^[���   ;��z�����]�������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u������EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;��ӌ����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��@���_^[���   ;��0�����]� ����������������������������������������������U����   SVWQ������<   ������Y�M�h�   �������E�}� t�E샸�    u�M�0����E�9��E�P�����Q�U싂�   �Ѓ�;�舋��P�M��������������E_^[���   ;��a�����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u������E�P�M싑�   �҃�;��Ǌ��_^[���   ;�跊����]����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u���EP�M�Q�U싂�   �Ѓ�;��&���_^[���   ;�������]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��|���_^[���   ;��l�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��Ј��_^[���   ;��������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��(���_^[���   ;�������]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3��+��EP�MQ�UR�EP�M�Q�U싂�   �Ѓ�;��x���_^[���   ;��h�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u����#��EP�MQ�U�R�E싈�   �у�;��φ��_^[���   ;�迆����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;�� ���_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��l���_^[���   ;��\�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;�輄��_^[���   ;�謄����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u������EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��x���_^[���   ;��h�����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��؂��_^[���   ;��Ȃ����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��8���_^[���   ;��(�����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;�蘁��_^[���   ;�舁����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;�����_^[���   ;��܀����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��H���_^[���   ;��8�����]�����������������������������������������U����   SVWQ������>   ������Y�M�h�   �������E�}� t�E샸�    u�M������E�N��EP�M�Q�����R�E싈�   �у�;�����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��\����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u�#��EP�MQ�U�R�E싈�   �у�;��~��_^[���   ;��~����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��~��_^[���   ;��~����]�����������������������������������������U����   SVWQ������>   ������Y�M�h�   �c������E�}� t�E샸�    u�M�̀���E�N��EP�M�Q�����R�E싈�   �у�;��d}���U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��,}����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u�#��EP�MQ�U�R�E싈�   �у�;��|��_^[���   ;��r|����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�P�M싑�   �҃�;���{��_^[���   ;���{����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��D{��_^[���   ;��4{����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u���#��EP�MQ�U�R�E싈�   �у�;��z��_^[���   ;��z����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u�,����E�$�EP�MQ�U�R�E싈�   �у�;���y��_^[���   ;���y����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��@y��_^[���   ;��0y����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��x��_^[���   ;��x����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h   ��������E�}� t�E샸    u3����EP�M�Q�U싂   �Ѓ�;���w��_^[���   ;���w����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h  �C������E�}� t�E샸   u3����E�P�M싑  �҃�;��Xw��_^[���   ;��Hw����]�����������������������������������������U����   SVWQ������>   ������Y�M�h  �������E�}� t�E샸   u�����$�M�Ak���E�J��E�P�����Q�U싂  �Ѓ�;��v���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��hv����]� ������������������������������������������������������U����   SVWQ������>   ������Y�M�h  �������E�}� t�E샸   u�����$�M�Qj���E�J��E�P�����Q�U싂  �Ѓ�;��u���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��xu����]� ������������������������������������������������������U����   SVWQ������>   ������Y�M�h  ��������E�}� t�E샸   u�����$�M�ai���E�J��E�P�����Q�U싂  �Ѓ�;���t���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��t����]� ������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h  ��������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;���s��_^[���   ;���s����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h  �3������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;��Fs��_^[���   ;��6s����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h  �������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;��r��_^[���   ;��r����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h   ��������E�}� t�E샸    u3����E�P�M싑   �҃�;��r��_^[���   ;���q����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h$  �S������E�}� t�E샸$   u3����EP�M�Q�U싂$  �Ѓ�;��dq��_^[���   ;��Tq����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h(  �������E�}� t�E샸(   u3��'��EP�MQ�UR�E�P�M싑(  �҃�;��p��_^[���   ;��p����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h,  �������E�}� t�E샸,   u�'��EP�MQ�UR�E�P�M싑,  �҃�;��p��_^[���   ;���o����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h0  �S������E�}� t�E샸0   u3����E�P�M싑0  �҃�;��ho��_^[���   ;��Xo����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h4  �������E�}� t�E샸4   u3����EP�M�Q�U싂4  �Ѓ�;���n��_^[���   ;��n����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h8  �������E�}� t�E샸8   u3��#��EP�MQ�U�R�E싈8  �у�;�� n��_^[���   ;��n����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h<  �c������E�}� t�E샸<   u�'��EP�MQ�UR�E�P�M싑<  �҃�;��nm��_^[���   ;��^m����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h@  �������E�}� t�E샸@   u�'��EP�MQ�UR�E�P�M싑@  �҃�;��l��_^[���   ;��l����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�hD  �������E�}� t�E샸D   u3����E�P�M싑D  �҃�;��l��_^[���   ;��l����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�hH  �c������E�}� t�E샸H   u3����EP�M�Q�U싂H  �Ѓ�;��tk��_^[���   ;��dk����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�hL  ��������E�}� t�E샸L   u3��#��EP�MQ�U�R�E싈L  �у�;���j��_^[���   ;���j����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�hP  �������E�}� t�E샸P   u3��'��EP�MQ�UR�E�P�M싑P  �҃�;��j��_^[���   ;��j����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�hT  �c������E�}� t�E샸T   u���'��EP�MQ�UR�E�P�M싑T  �҃�;��li��_^[���   ;��\i����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�hX  �������E�}� t�E샸X   u�0����E�$�EP�MQ�UR�E�P�M싑X  �҃�;��h��_^[���   ;��h����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j<�������E�}� t	�E�x< u� ��EP�MQ�U�R�E�H<�у�;��h��_^[���   ;��h����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M�j@�f������E�}� t	�E�x@ u3����EP�M�Q�U�B@�Ѓ�;��}g��_^[���   ;��mg����]� �������������������������������������������U����   SVW��4����3   ������j�K   ���E��}� u3���E���H��;���f��_^[���   ;���f����]�����������������������U����   SVW��@����0   ������h�/�EPh�� ��x����_^[���   ;��f����]�������������������������U����   SVW��(����6   ������E�8 u�>j�q������E��}� u�)�E��M��E�P�M��Q�҃�;��f���E�     R��P�|6�Q��XZ_^[���   ;���e����]Ð   �6����   �6i ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3��$��EP�MQ�UR�EP�U�M��B��;��5e��_^[���   ;��%e����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u���EP�MQ�U�M��B��;��d��_^[���   ;��d����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j�v������E�}� t	�E�x u���EP�MQ�U�M��B��;��d��_^[���   ;���c����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3��,��EP�MQ�UR�EP�MQ�UR�E�M��P��;��mc��_^[���   ;��]c����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �6������E�}� t	�E�x  u3��(��EP�MQ�UR�EP�MQ�U�M��B ��;���b��_^[���   ;��b����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u3��$��EP�MQ�UR�EP�U�M��B$��;��b��_^[���   ;��b����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3��$��EP�MQ�UR�EP�U�M��B(��;��ua��_^[���   ;��ea����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�F������E�}� t	�E�x, u3��6��E$P���E�$���E�$�MQ�UR�EP�U�M��B,��;���`��_^[���   ;��`����]�  �������������������������������������������������U����   SVWQ��(����6   ������Y�M�j0�������E�}� t	�E�x0 u3��(��EP�MQ�UR�EP�MQ�U�M��B0��;��`��_^[���   ;��`����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4��������E�}� t	�E�x4 u3��9��E(P���E �$�MQ�UR�EP�MQ�UR�EP�U�M��B4��;��P_��_^[���   ;��@_����]�$ ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u�����EP�MQ�U�M��B8��;��^��_^[���   ;��^����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�v������E�}� t	�E�x< u���EP�MQ�U�M��B<��;��^��_^[���   ;���]����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j@��������E�}� t	�E�x@ u3����EP�MQ�U�M��B@��;��}]��_^[���   ;��m]����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jH�F������E�}� t	�E�xH u3����EP�MQ�U�M��BH��;���\��_^[���   ;���\����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jD�������E�}� t	�E�xD u3����EP�MQ�U�M��BD��;��=\��_^[���   ;��-\����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jL�������E�}� t	�E�xL u���!��EP���E�$�U�M��BL��;��[��_^[���   ;��[����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jP�f������E�}� t	�E�xP u3����EP�MQ�U�M��BP��;���Z��_^[���   ;���Z����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jT��������E�}� t	�E�xT u3��$��EP�MQ�UR�EP�U�M��BT��;��UZ��_^[���   ;��EZ����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�jX�&������E�}� t	�E�xX u3��,��EP�MQ�UR�EP�MQ�UR�E�M��PX��;��Y��_^[���   ;��Y����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u3��,��EP�MQ�UR�EP�MQ�UR�E�M��P\��;���X��_^[���   ;���X����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u�Zf���M��A�E��x u3���E�P�MQ�UR�EP�M��I��E��_^[���   ;��MX����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�EP�MQ�U��J�M���E���P�?X����_^[���   ;��W����]� ����������������������������U����   SVWQ��4����3   ������Y�M��E��x u�:e���M��A�E��x t�EP�MQ�U��J�=��_^[���   ;��9W����]� ���������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t+�MQ�UR�EP�MQ�UR�EP�M��I�_����0����
ǅ0���    ��0���_^[���   ;��V����]� �����������������������������������U����   SVWQ��0����4   ������Y�M��E��x t'�MQ�UR�EP�MQ�UR�E��H�_����0����
ǅ0���    ��0���_^[���   ;���U����]� ���������������������������������������U����   SVWQ��0����4   ������Y�M��E��x u�jc���M��A�EP�MQ�UR�EP�M��H����u3��<�E��x t#�MQ�UR�EP�MQ�U��J�T����0����
ǅ0���    ��0���_^[���   ;��)U����]� �������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t#�MQ�UR�EP�MQ�U��J�\R����0����
ǅ0���    ��0���_^[���   ;��}T����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t5�M$Q���E�$���E�$�UR�EP�MQ�U��J�`F����0����
ǅ0���    ��0���_^[���   ;���S����]�  �����������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t'�MQ�UR�EP�MQ�UR�E��H��O����0����
ǅ0���    ��0���_^[���   ;��)S����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� 8�M���7��_^[���   ;��R����]�������������������������U����   SVWQ��4����3   ������Y�M��M��K���E��t�E�P�L>�����E�_^[���   ;��JR����]� ������������������������U����   SVWQ��(����6   ������Y�M��M�7���E�M��Q�P�E�M��Q�P�E�    �	�E���E�E��M�;H}�E��H�U��P�M�@����u3���͸   _^[���   ;��Q����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��} |$�E��M;H}�} |�E��M;H}�E;Eu�"�E��H�U��P�M��Q�E��Q��9����_^[���   ;���P����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E;E}	�E���E�} |$�E��M;H}�} |�E��M;H}�E;Eu�/�E��H�U���E�EP�M��<<����t�EP�M�Q�M���c��_^[���   ;��P����]� �������������������������������������������U����   SVWQ������9   ������Y�M��E��x u�E��H�M��%�E��x t�E��H�U�J�M���E��H��M��}� u3��]��h@����P�M���Q�U��BP��*�Q��  �Ѓ�;��MO���E�}� u3���E��M�H�E��M��H�   _^[���   ;��O����]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��P;Qu�M��E����u3��&�E��H�U��B�U���E��H���U��J�   _^[���   ;��eN����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��M;H}�EP�MQ�M��J���#�E��H;M}j �M���<����EP�M��<��_^[���   ;���M����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3���E��H�U�E���   _^[��]� ���������������������������U����   SVWQ��(����6   ������Y�M��E��M;H~	�E��H�M�} }�E    �E��M��P;Qu�M��C����u3��Z�E��H�M��	�E���E�E�;E~�E��H�U��B�U�u�L�����ԋE��H�U�E���E��H���U��J�   _^[���   ;��`L����]� ��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3��E�E��H���U��J�	�E���E�E��M;H}�E��H�U��B�U�u�L����Ѹ   _^[��]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��<8��P�M��/7��_^[���   ;��$K����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E��M�;H}�E��H�U��;Eu�E���ԃ��_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E���P�A�����E��@    �E��@    �M��A    _^[���   ;��J����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��@    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M��E��H��Q�M���[���E�}� t�E��H��Q�M��W5���E�_^[���   ;��II����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H}�E��H�U���3�_^[��]� �������������������U����   SVWQ��$����7   ������Y�M��EP�M���Y��j�E��HQ�U��BP�M���-��R��P� T�4��XZ_^[���   ;��dH����]� ��   T����   Tsort ���������������������������������������U����   SVWQ��4����3   ������Y�M��M���\���E�� ��E��M�H�E�_^[���   ;���G����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�Ѓ�;��mG��_^[���   ;��]G����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�� ��E�_^[��]���������������������������U����   SVWQ��$����7   ������Y�M��EP�M���W��j�E��HQ�U��BP�MQ�M��Q��R��P��U�82��XZ_^[���   ;��F����]� ��   �U����   �Usort �����������������������������������U����   SVWQ��4����3   ������Y�M��E�� ��M����O���M����O���E��@    �M���5���E�_^[���   ;���E����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E�� ��E��@    �E��@    �E�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��M���R���E��t�E�P��0�����E�_^[���   ;���D����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��7Z���E��t�E�P�0�����E�_^[���   ;��D����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� ��M��K���M�����Q���M�����Q��_^[���   ;��D����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E����M��A�E����M��A�E��@    _^[��]���������������������������U���   SVWQ�� ����@   ������Y�M��M��L���E��}� tm�M��R���E�}� tM�E��������������������� t%��j��������������;���B���� ����
ǅ ���    �E�    �E�E�덋M���2��_^[��   ;���B����]����������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t�M��Q�z t�E��H��0����
ǅ0���    ��0���_^[��]������������������������������������U����   SVWQ��0����4   ������Y�M��E����M�9At�U��B��0����
ǅ0���    ��0���_^[��]���������������������������U����   SVWQ������9   ������Y�M��M��J���E��}� t�M��P���E�M��H���E�E���_^[���   ;��=A����]������������������������������U����   SVWQ������:   ������Y�M��E�    �M��J���E��}� tD�E�M�U���U�;�uǅ���   �
ǅ���    ����� t�E���M���O���E��3�_^[���   ;��@����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E�M��Q�P�E����M�A�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E����M�A�E�M��Q�P�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ������9   ������Y�M��E�    �M��XH���E���M��hN���E��}� t�E���E���E�_^[���   ;���>����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� ��M���E��_^[���   ;��>����]�������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E�H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t;�E��x t2�E��H�U��B�A�E��H�U��B�A�E��@    �M��A    _^[��]�����������������������������������U����   SVW��4����3   ������E��M��E�M���E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M�jh�  �M�_7���EP�MQ�M���4��_^[���   ;��:<����]� ������������������������U����   SVWQ��(����6   ������Y�M��E����M��BX��;���;��P�M�6+����t$ǅ,���   ��,���P�MQ�|+�����   ��EP�MQ�UR�EP�M��5��_^[���   ;��;����]� ����������������������������������������U����   SVW��@����0   ������E�M��E��E_^[��]��������������������������U����   SVWQ��0����4   ������Y�M�j �M�v:��� ��0�����0����  t�7�5�3�E��x u*j h�  �M�7����uj h�  �M�7����t3�� �EP�MQ�UR�EP�MQ�UR�M��q@��_^[���   ;��b:����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �EP�N2����_^[���   ;���9����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��@   �   _^[��]� ���������������������U����   SVWQ��4����3   ������Y�M��E��@   _^[��]� ��������������������������U���`  SVWQ�������X   ������Y�M��}`��u
�E��@   �}��   �E�E�j �M��c8���8�  u)�<H��P�M��<:��jh�  �M�3���   �  �vj �M��(8���8�  u*��EP�MQ�U���M��P��;��k8���   �j  �:j �M���7���8�  tj �M���7���8ujh�  �M�43���E��@    �}�  �E�E��E��H���U��Jj	�E����M��BX��;���7��P�G�����E��E�    �}� tj �M��k=���EȋE��M�;H��  �E��x ��  j h�  �M�4����uj h�  �M�o4�����s  j h�  �M�x2���}� tj �M��=���EȋE��MȉH�M��=���} t�M��nK����uǅ����   �M������������)  �EP�*.�����M���K��j�M��/K��P�M�1����t�����K���E��|����M��
K���E��E��t����E�   �M��B��������������t������t������t��E�   ��E�   ��E�   ��E�    ��%����t��� t��t����M����t���P�M����M��BX��;��G6��P�L!������t��� t��t����_����t����(<���M�� <���M������EP�MQ�UR�EP�M��8��R��P��f�!��XZ_^[��`  ;���5����]�    �f����   �f����   �ft���   �fmd mu pActive ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q��*�BH���  �у�;��d4��_^[���   ;��T4����]� ����������������������������������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M���:���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��3����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;���2����}�EP�M�Q�U�R�M��:�����U��������_^[��,  ;��2����]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M��J���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��z0����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��J0����}�E�P�M�Q�U�R�M��u�����U��������_^[��8  ;��0����]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M��}���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;���-����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��-����}�E�P�M�Q�U�R�M�������U��������_^[��8  ;��c-����]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��u�EP�MQ�UR�M������83��} ����t�EP�MQ�UR�M�������EP�MQ�UR�M��/��_^[���   ;���+����]� �������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  �Ek� E�E���E�P�MQ�U���M����;��!+���Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;��*���Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��n*����t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;��&*����]� ����������������������������������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u�E� ����3���  �Ek� E�E���E�P�MQ�U���M����;��H)���Eȃ}� u
�E��  ��}� }�E�     3��  �E�   �E���E��E�    �E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;���(���Eȃ}� uS�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��(����t�
��E��E�뷋E���   ��}� }�Eԃ��E��	�Eԃ��E��D����}� ~�Eԃ��M���E�Mԉ�E�;M}F�E�M�M�M���E�P�MQ�U���M����;���'����|h��4��9P������E�8 ~I�E����MM�M���E�P�MQ�U���M����;��'����h��4��?P�F����3�_^[��  ;��~'����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M����_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��M�2,���E_^[���   ;��%����]� ����������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]�  ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��(����6   ������Y�M��} u3��]��EP�M���M��B@��;���#���E�}� u3��6�M�������P�EP�MQ��*�B0���   �у�;��#���M�����_^[���   ;��#����]� ������������������������������������������������U����   SVWQ������=   ������Y�M���EP��*�Q0�B�Ѓ�;��+#���E�}� tM�E쉅 ����� ������������� t%��j��������������;���"��������
ǅ���    �E�    _^[���   ;��"����]� ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�j�E�Q�G������t�   �3�_^[���   ;��� ����]� ��������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�j�E�Q�[������t�   �3�_^[���   ;�������]� ��������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVW��@����0   �������EP�MQ��*�B���  �у�;����_^[���   ;��	����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP��*�Q���  �Ѓ�;����_^[���   ;������]����������������������������������U����  SVW��(����v   ������ǅ ���    �}( uǅ0���    �M�1����0����!  �E�    �M��(������  �M������M��+������   �EP��H�����2���� ���j h����������'���� ���P��l����2���� ���j j���H���Q��l���R������P�c3������ ���P������Q������� ���P������R�p������ ��� P�M��=���������uǅ(���   �
ǅ(���    ��(�����?����� ����� t�� ���ߍ������_
���� �����t�� ��������B
���� �����t�� �����������%
���� �����t�� ������l����
���� �����t�� �����������0���� �����t�� ������H�����	����?�����t(�E(P�M$Q�M����P�UR�EP�MQ�������E��M��(���!�E(P�M$Qj �UR�EP�MQ�������E��E�������M�/�������R��P������XZ_^[���  ;�������]ÍI    ������   ��icon �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������EP�MQj �UR�EP�MQ�����_^[���   ;�������]���������������������������������U���  SVW��H����n   ������} u3��g  j h�   ��<���P�c������$���P�M��M�B��;��>����$�����$����t9j ��$���P�MQ���������u ǅL���    ��$����-����L�����   �E��\����E��|����E�E��E��<���ǅ@������E�L��E�_��E�k��E����E�ݝ�E�K��E�׀�E���E�Q��E�ϡ�E�(��E�u��E����E�B��E���E����E�G��E�p��E�d��EЏ�h�   ��<���P�MQ�URj	�]������X�����$����,����X���R��P�x����XZ_^[�ĸ  ;�������]Ð   ��<����   ��$���   ��description np �������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q��*�B���   �у�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$���E�$�MQ�U�R��*�H���   �҃�;��O��_^[���   ;��?����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q���   �Ѓ�;�����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P��*�Q���   �Ѓ�;��X��_^[���   ;��H����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P��*�Q���   �Ѓ�;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���   �҃�;��a��_^[���   ;��Q����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP��*�Q�Bp�Ѓ�;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���  �҃�;��q��_^[���   ;��a����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���  �҃�;��q��_^[���   ;��a����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R��*�H���  �҃�;�����_^[���   ;�������]� ������������������������������̋�`<����������̋�`L����������̋�`����������̋�` ����������̋�`0����������̋�`P����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`����������̋�`����������̋�`,�����������u�U��� PRSVW�Ej P�>����_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR�!�����E�@���E�;|�_^[��]���������������������������̋�U��V���t!��tS�]��tW�̋�����F�V�3_[^]� �������������̋�U��QSVW��3���;�tR�}�9>~K��    �F�8�����9T�u�D8�9t�N�T�ERP�a��������̋E�@���E�;|������̋u3��ƅ�tV�@G��u���tJ9u9Vu
9Vu9Vt�MWVQ�T��������̋F9T0�t�MWVQ�8��������̋vO��u�_^[��]� �����������������������������������������������������������̀=�/ uj jj j j ��/����P������������������������������jjj j j ������������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������������̋�U��Q�M��EP�M�Q��������]� ����������������̋�U��Q�M��E�� �M�Q���������]��������������̋�U��Q�M��M�������E��t�M�Q��������E���]� �����������������̋�U��Q�M��EP�M�Q�.�������]� ����������������̋�U��Q�M��E�P�B������]�������̋�U��Q�M��E���	P�M��	Q��������������]� �������������������̋�U��Q�M��E���	P�M��	Q����������؋�]� ��������������������̋�U��Q�M��E���	P�M��	Q�`�����3҅���]� �����������������̋�U��Q�M��E�����]�������������̋�U��Q�M��E�� �E���]� ��������������������̋�U��Q�M��E���]� �������������̋�U���g���} t�0�����]�������̋�U����F���$������S������F���P���i�������ң]�������������������������������������̋�U��Q��/�E��M��/�E���]������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �}��   ������u3��  �����u����3��  ������a� U�K����/�	����}��������3��i  �����|�����|j �������t��������T���3��3  j�n������/����/�  �} um�=�/ ~X��/����/�E�    �=40 u����Y����-��������E������   ��} u�=��t�����3��   �   �}��   �����h�   h(jh  j������E�}� tV�U�R��P��/Q��a�Ѕ�t%j �U�R�&������a�M��U��B�����j�E�P������3���3����}u
j ��������   �M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��}u�����EP�MQ�UR�   ��]� �����������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e��E�   �} u�=�/ u3��N  �E�    �}t�}uT�=$ t�EP�MQ�UR�$�E�}� t�EP�MQ�UR�m���E�}� u�E�    �E������E���   �EP�MQ�UR����E�}u=�}� u7�EPj �MQ�����URj �EP����=$ t�MQj �UR�$�} t�}u@�EP�MQ�UR������u�E�    �}� t�=$ t�EP�MQ�UR�$�E��E������8�E���U��E�P�M�Q������Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    ����E�    �EP�Y   ���E��E������   ��_��ËE�M�d�    Y_^[��]������������������������������������������̋�U����UP��a�E��UQ��a�E��U�;U�r�E�+E�����s3���   j�M�Q�F������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}hdj�E�P�M�Q�������E��}� u:�U���U�E�;E�r%h�   hdj�M�Q�U�R������E��}� u3��Q�E�+E����M����U��E��E��M�Q��a�U�UR��a�M���U����U��E�P��a�U�E��]�����������������������������������������������������������������������������������������������̋�U��EP����������؃�]��������������������̋�U��Qh�   hdjjj ������E��E�P��a�U�U�U�}� u�   ��U��    3���]�������������������������;hu���1�������������������̃=�S ��
�����\$�D$%�  =�  u�<$f�$f��f���d$��
��� �~D$f(�f(�f(�fs�4f~�fT�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�������D$��~D$f��f(�f��=�  |!=2  �fT��\�f�L$�D$����f��fV�fT�f�\$�D$�������������������������������������������������������������������������������̃=�S t-U�������$�,$�Ã=�S t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������������������������������������������������������̋T$�L$��ti3��D$��u���   r�=�S t�e���W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̋�U��Qj j j�X5P�MQ�� �����E��E���]������������������������̋�U��j�EP�x�����]������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̋�U������]�h��  h?  ��������E��E%�  =�  ��   ���E�$�o������E�}�t�}�t!�}�t3�Jh��  �M�Q�������E�   h��  �U�R�������E���i�E�P���E�$j�D������P�M�Q�E������$���E�$jj�7������&�U������U�E�E�h��  �M�Q�������E���]��������������������������������������������������������������������̺ ����� �.	�����������z�����������������̋�U��Q��<P��a�E��}� t�U�j������jj �U������$����]�������������������̋�U��Q�E�    ��<P��a�E��MQ��a��<�E���]��������������̋�U���<P��a]�������������̋�U��E��w$��p���
���tRP�EQP�D   ��]ú�R�   P�E�   QP�$   ��]�������������������������������̋�U���@  �h3ŉE��ES�]VW�}S������������ǅ����    �g������������uS�
�����������5�aj j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ����h  ��  ����������t%���������
PSQW�}  �����"  2��������� ������u���  ��t��a����   h  ������R������Ph  ������Q���S��������t-������������RWh�������P�EQ������RP���   �=�aj j h
  ������Qj�������Rj h��  ���ׅ�t������j j h
  ������Pj�������Qj h��  ���ׅ�t������������������������R�UPh`VQSR����������u̋M�_^3�[�l����]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h �h5�d�    P��$SVW�h1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@��a�	�   Ëe��E������E�M�d�    Y_^[��]��������������������������������������̋�U��j�h �h5�d�    P��$SVW�h1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@��a�	�   Ëe��E������E�M�d�    Y_^[��]����������������������������������������������������̋�U���  �h3ŉE��=x��E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ���
������A��u�Њ@��u�W������+�O�OG��u��������ȃ���
�Ȋ@��u�������+���O�OG��u������ȃ��_����x������SjPQ�������^[�M�3��a����]��������������������������������������������������������������������̋�U���D  �h3ŉE�S��V�uW�}�����������   h� b����   h�P��a��/����   ����   �M�Vh�Qh���$Rh��~ Wh�hH������h,Q�ЋV��$RW�E�P�M�Q��   ��8h(�U�Rh$�E�Ph������Q��a������R��/������������PjSQ������(_^[�M�3������]�h�jSW�������M�_^3�[������]�����������������������������������������������������������������������������̋�U����ESV�u�E��EW3�+ƉE����M��r�   ;�s&�0�U���Qh$R��/�E��E����GF�ɋM�E�y� � _^[��]���������������������������������̋�U���  �h3ŉE��=|��E��   SV����   �ȍq�A��u�+΃�:��   ww������3Ɋ�������A��u�Њ@��u�W������+�O�OG��u��������ȃ���Ȋ@��u�������+���O�OG��u������ȃ��_��,�|SjP�EP������^[�M�3��$����]�����������������������������������������������������������������������̸   ����������̋�U��E��w	��8]�3�]������̋�U��M��w�U��p��p]Ã��]�����������̋�U��M��/��/��/    ]�����������������̋�U��M��/��/��/    ]�����������������̡�/����������̡�/�����������u�U��� PRSVWh�h�jBhPj��������u�_^[ZX��]������������������������̋�U���]����̋�U��|�]����̋�U��j�h@�h5�d�    P���SVW�h1E�3�P�E�d�    j�D������E�    �E�x ��   ��/�M��E�/��U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�������/�M�M��U�z uh8j jXh�j��������u�랋M�QR�}������E�@    �E������   �j������ËM�d�    Y_^[��]������������������������������������������������������������������������̋�U��j�h`�h5�d�    P���SVW�h1E�3�P�E�d�    �E�x �L  h (  h	�hٰj �M��	Qj �������E�}� u3��   �U�R�������E��E��M����M���v�U�U���� u�M�M�� ��j�}������E�    �U�z ��   j�H������E܃}� ��   �E���P�,������E؋M�U؉Q�}� t[j h�   h�h(hp�E�P�M���Q�U�BP�o�����P��������M܋U�B��M܋U�B�A�M�U܉Q��E�P�������M�Q�������E������   �j�������ËU�B�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������̋�U��} u��EP�MQ�UR�EP�MQ����]������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    j�������E�    �E�x ��   ��/�M��E�/��U��U�}� tY�E�M�;Qu�E��M�Q�P�E�P�������2�M�M��U�z u!h8j h�   h�j���������u�뛋M�QR�f������E�@    �E������   �j������ËM�d�    Y_^[��]���������������������������������������������������������������������̋�U���E��u	� (  f�M�URh	�hٰ�EP�MQ�UR�;�����]���������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E�x �a  j��������E�    �M�y �*  h (  j �U��	Rj �������E�}� u"�E�    j��E�Phh��������E��  �M�Q�s������E��U��E����E���v�M�M���� u�E�E��  ��j� �����E܃}� ��   �E�    �M���Q�g �����E؃}� taj h4  h�h�h`�U�R�E���P�M�Q�s�����P��������U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P�!������M�Q�������E������   �j�������ËU�B�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    j��������E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P��������M�Q����������E������   �j������ËM�d�    Y_^[��]�����������������������������������������������̋�U��j jh�h�h(h   h   j �[�����P�������]�������������������������̋�U��j �EP�������]�����������̋�U����EP�M������M�R�J�������et�E���E�M�R���������u�E�Q��������xu	�U���U�E��M��M���������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M��������]������������������������������������������������̋�U��Q�M��E��@ �} ��   �����M��A�U��B�M��Pl��E��H�U��Ah�B�M��;�t�E��H�Qp#8u
�����M���U��B;8t�M��Q�Bp#8u������M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������������������������������������������������������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]�������������������̋�U��Q�M��E���]����������������̋�U��j �EP�,�����]�����������̋�U���V�EP�M������M���t*�E�0�M��v�������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M����������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M�����^��]�������������������������������������������������������������������̋�U��Q�E�������Az	�E�   ��E�    �E���]���������������������̋�U����} t$�EP�MQ�U�R�O������E�M���U��P��EP�MQ�U�R�\������E�M���]������������������������������̋�U��j �EP�MQ�UR�������]�������������������̋�U���D�h3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�������3Ƀ} ���Mă}� u!hj h�  h�j�q�������u̃}� u3�����    j h�  h�h|h�������   �  3�;E��ىM�u!hTj h�  h�j�	�������u̃}� u3�"����    j h�  h�h|hT�A������   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�������Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3��a�����]��������������������������������������������������������������������������������������������������������������������̋�U���@�E�    �E P�M�����3Ƀ} ���M܃}� u!hj h3  h�j�g�������u̃}� u@�����    j h3  h�h�h�������E�   �M��.����E���  3�;E��ىM�u!hTj h4  h�j���������u̃}� u@�����    j h4  h�h�hT�*������E�   �M������E��}  3��} ����#E��	;E��ىM�u!hj h<  h�j�m�������u̃}� u@����� "   j h<  h�h�h�������E�"   �M��4����E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�V  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��G�������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  h�h�h@h8�U�R�E�P�������P�h������M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE����?��t �U����0uj�M��Q�U�R�������E�    �M��7����Eċ�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M������} }�E    3Ƀ} ���M��}� u!hj h�  h�j�c�������u̃}� u@�|����    j h�  h�h$h�������E�   �M��*����E���  3�;E��ىM�u!hTj h�  h�j���������u̃}� u@�����    j h�  h�h$hT�&������E�   �M������E��g  �E�  �M��;M��ډU�u!h�j h�  h�j�o�������u̃}� u@����� "   j h�  h�h$h��������E�"   �M��6����E���  �M��Q�4����%�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ��������E��}� t�U� �E��E��M������E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ�:������E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M������E���  �M��Q�?�������� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4����%�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M��_�������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U������E�U��E܅���   �} ~}�M��Q���� #E�#U��M������f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U������E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M��G���f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4�X���%�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�s�������0�M��U���Uj h�  �E�P�M�Q�#����E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�����Ѓ�0�E��M���Mj jd�U�R�E�P������E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P������ȃ�0�U�
�E���Ej j
�M�Q�U�R�����E��U��E���0�M��U���U�E�  �E�    �M��I����E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ������]���������̋�U��j �EP�MQ�UR�EP�MQ�>�����]�����������̋�U���D�h3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�������3Ƀ} ���Mă}� u!hj h*  h�j聽������u̃}� u3�����    j h*  h�h<h�������   ��   3�;E��ىM�u!hTj h+  h�j��������u̃}� u3�2����    j h+  h�h<hT�Q������   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP��������Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�   ���EȋEȋM�3�������]�����������������������������������������������������������������������������������������������������������̋�U���4�E�H���M��UR�M������3��} ���E�}� u!hj h�  h�j蒻������u̃}� u@�����    j h�  h�hTh��������E�   �M��Y����E��  3�;U��؉E�u!hTj h�  h�j��������u̃}� u@�6����    j h�  h�hThT�U������E�   �M�������E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P��  ���M��0�U����U���E�M�H�M��} ��   j�U�R�  ���M�赹��� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�  ���EPj0�M�Q�������E�    �M������EЋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U���P�h3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P������3Ƀ} ���M��}� u!hj ho  h�j�M�������u̃}� u3�f����    j ho  h�hlh�������   �i  3�;E��ىM�u!hTj hp  h�j��������u̃}� u3������    j hp  h�hlhT�������   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�������E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�?������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ��������M�3��������]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�������]�����������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�������E��{�}fu!�E P�MQ�UR�EP�MQ�o������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ耯�����E��#�U R�EP�MQ�UR�EP�MQ�"������E��E���]������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�����������������������̋�U��} t#�EP蘸������P�MQ�UUR�������]����������������̋�U��Q�E�    �	�E����E��}�
s�M����R��a�M�����ԋ�]�����������������̋�U��j ��a]�����������������̋�U���b]� ����������������̋�U��EP��Q�b��]� �������������������̋�U�졸]����̋�U��Q��P�b�E��}� u ��/Q��a�E��U�R��P�b�E���]������������������������������̋�U��EP�MQ��/R��a��]� ���������������̋�U���h��b�E��}� u����3���  h��E�P��a��/h��M�Q��a��/h��U�R��a��/h��E�P��a��/�=�/ t�=�/ t�=�/ t	�=�/ u,��/���b��/�b��/�b��/�b���=��t��/Q��R�b��u3���   �ӷ����/P��a��/��/Q��a��/��/R��a��/��/P��a��/������u�m���3��   h����/Q��a�У��=��u	�?���3��rh  h�jh  j�i������E��}� t�U�R��P��/Q��a�Ѕ�u	�����3��(j �U�R�p�������a�M���U��B�����   ��]������������������������������������������������������������������������������������������������������������������������������������̋�U��=��t��P��/Q��a���������=��t��R�b�������v���]����������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    h��b�E�E�@\p1�M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@hj谰�����E�    �M�QhR�b�E������   �j�������j�y������E�   �E�M�Hl�U�zl u�E���Hl�U�BlP�������E������   �j�`�����ËM�d�    Y_^[��]��������������������������������������������������������������������������̋�U���� b�E���P�D����ЉE��}� u}j h�  h�jh  j�c������E��}� tW�M�Q��R��/P��a�Ѕ�t%j �M�Q�v�������a�U���E��@�����j�M�Q�.������E�    �U�R�b�E���]�����������������������������������������������������������̋�U��Q�����E��}� u
j��������E���]�����������̋�U��j�h�h5�d�    P���SVW�h1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P�O������M܃y, tj�U܋B,P�5������M܃y4 tj�U܋B4P�������M܃y< tj�U܋B<P�������M܃y@ tj�U܋B@P��������M܃yD tj�U܋BDP��������M܃yH tj�U܋BHP�������M܁y\p1tj�U܋B\P������j葭�����E�    �M܋Qh�U��}� t%�E�P�$b��u�}�tj�M�Q�Q������E������   �j�q������j�3������E�   �U܋Bl�E�}� t4�M�Q�������U�;�t�}��t�E�8 u�M�Q�b������E������   �j�������j�U�R�������M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��=��tO�} u)��P�b��t��Q��R�b�ЉEj ��P��/Q��a�ЋUR�ӻ���=��tj ��P�b]������������������������������������������̋�U����a]���̋�U���(b]���̋�U��Q�EP�MQ�UR�X5P�MQ�r������E��E���]������������������̋�U��j j j�EP�MQ�;�����]�������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�D   ���E��}� u�}� t������t
�����M���E���]������������������������̋�U��Q�EP�MQ�UR�EP�MQ�   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP�O�������u�} t	�M�   3��뗋�]�����������������������������̋�U��j j j�EP�4�����]�������̋�U��j�h@�h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    j膩�����E�    �=�/ vU��/��9�/u6������u!h�j h  h(j��������u���/    ���/����/���E؃=��t�M�;�u̃=�  tu�UR�EP�M�Q�UR�EPj j�� ����uP�} t%�MQ�URh�j j j j �	�������u�� h�h� j j j j ��������u��D  �U����  ��t����u�E�   �}�v3�MQh�j j j j螧������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t hTh� j j j j�B�������u̋M��$�MԋU�R�������E܃}� u�} t	�E�    �r  �������}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+�/;Mv��/U��/�
��/������/E��/��/;�/v��/��/�=�/ t��/�M܉H�	�U܉�/�E܋�/��U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉�/j��R�E܃�P�S�����j��Q�U�E܍L Q�6������UR��P�M܃� Q�������U܃� �U��E������   �j�]�����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�(������E��}� u�}� t�������t
������U���E���]����������������������������̋�U��Q�} v�����3��u;Es�����    3��K�E�E�E�MQ�UR�EP�MQ�X5R�EP��������E��}� t�MQj �U�R�������E���]���������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR踤�����E��}� u�}� t�������t
�����M���E���]������������������������̋�U��Qj j j�EP�MQ�UR�؛�����E��E���]����������������������̋�U��j�h`�h5�d�    P���SVW�h1E�3�P�E�d�    j�$������E�    j�EP�MQ�UR�EP�MQ�b   ���E��E������   �j������ËE�M�d�    Y_^[��]����������������������������������������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R譜�����  �} t�}� u�EP�MQ�E�����3��  �=�/ vV��/��9�/u6�i�����u!h�j h�  h(j�Ԡ������u���/    ���/����/���U�=��t�E�;�u̃=�  ty�MQ�UR�E�P�MQ�U�R�EPj�� ����uR�} t%�MQ�URh<j j j j �ɠ������u�� hh� j j j j 觠������u�3��  �}��v`�} t)�UR�EP�M�Qh�j j j j�m����� ��u���E�Ph�j j j j�L�������u�������    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh`j j j j��������u�� hTh� j j j j�Ο������u��Qj��R�E�����P�  ����t1�MQh j j j j荟������u��%����    3��t  �EP��������u!h�j h  h(j�Þ������u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h j h#  h(j�n�������u��d�M�Q����  ��u�E%��  ��u�E   �M��/;Qs1�EPh�j j j j衞������u��9����    3��  �} t%�U���$R�E�P�͠�����E��}� u3��_  �#�M���$Q�U�R�_������E��}� u3��:  3�u��������}� u|�=�/�s9�U��/+B��/���+�/;M�v��/U���/�
��/�����E���/+H��/��/U���/��/;�/v��/��/�U��� �U�E��M�;Hv$�U��E�+BP��Q�U��E�BP�������j��Q�U�U�R��������}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!hHj h�  h(j�u�������u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8��/;M�t!hj h�  h(j��������u̋E��H��/�U��z t�E��H�U����7��/;M�t!h�j h�  h(j�˛������u̋E����/�=�/ t��/�E��B�	�M���/�U��/��M��A    �U���/�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es�����    3��g�E�E�E��} t�MQ�[������E��UR�EP�MQ�U�R�EP� ������E�}� t �M�;M�s�U�+U�Rj �E�E�P�K������E��]����������������������������������������������������̋�U��Qj j j�EP�MQ�߶�����E��E���]����������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E��}� u!h�j h�  h(j耘������u̃}� u-虻���    j h�  h(h�h�踲����3��c�}�v�f����    3��Nj�Y������E�    j �UR�EP�MQ�UR�EP�������E��E������   �j�L�����ËE�M�d�    Y_^[��]�������������������������������������������������������������������̋�U��j�EP������]�����������̋�U��j�h��h5�d�    P��SVW�h1E�3�P�E�d�    j�d������E�    �EP�MQ蒣�����E������   �j�h�����ËM�d�    Y_^[��]����������������������������������̋�U��Q�=�/ vU��/��9�/u6�!�����u!h�j h  h(j茖������u���/    ���/����/�} u�l  �}uOj��P�M�����Q�	  ����t/�URhp"j j j j訖������u��@����    �  �=�  tDj j j �MQj �URj�� ����u%hP"h� j j j j �P�������u���  �MQ��������u!h�j h*  h(j蓕������u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!h�!j h0  h(j�5�������u̋����m  j��P�M���Q�k  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��<Ph !j j j j�8�����(��u��<�U��� R�E��HQ�U��B%��  ��<Qhx j j j j������� ��u�j��P�M��Q�E��L Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��<Ph�j j j j�~�����(��u��<�U��� R�E��HQ�U��B%��  ��<Qhj j j j�@����� ��u̋E��xue�M��y����u	�U��z t!hxj hi  h(j�z�������u̋M��Q��$R��P�M�Q�W������U�R�צ�����Q  �E��xu�}u�E   �M��Q;Ut!h0j hw  h(j�	�������u̋M���/+Q��/������   �M��9 t�U���M��Q�P�6��/;E�t!h�j h�  h(j覒������u̋U��B��/�M��y t�U��B�M����5��/;E�t!h�j h�  h(j�X�������u̋U����/�M��Q��$R��P�M�Q�+������U�R諥�����(�E��@    �M��QR��P�M��� Q���������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�EP�E�����]�����������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E܃}� u!h�j h�  h(j�0�������u̃}� u1�I����    j h�  h(h�"h��h���������8  �=�/ vV��/��9�/u6�J�����u!h�j h�  h(j赏������u���/    ���/����/j軐�����E�    �UR觑������u!h�j h�  h(j�X�������u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!h�!j h�  h(j���������u̋E��xu�}u�E   �M��Q�U��E������   �j�#�����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������̋�U��Q���E��M���E���]������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    j�������E�    �EP���������te�M�� �M�U�B%��  ��tC�M�yt:�U�B%��  ��t*�M�yt!h�!j h?  h(j�V�������u̋E�M�H�E������   �j蓡����ËM�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�� �E��M�� �E���]������������������̋�U��� ]����̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�����������������������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    ����u
�   ��  j�0������E�    �Ŏ���E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$�x�h�%h� j j j j �&�������u��   h`%h� j j j j ��������u��dh8%h� j j j j �ߋ������u��Bh%h� j j j j 轋������u�� h�$h� j j j j 蛋������u��E�    ��  �E�   ��/�E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��<�U���E��$j��P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh !j j j j 豊����(��u��-�E�� P�M�QR�E�Phx j j j j 肊���� ��u��E�    j��R�E�H�U�D
 P�2�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph�j j j j ������(��u��-�U�� R�E�HQ�U�Rhj j j j ������ ��u��E�    �M�y ��   �U�BP��Q�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� Rh$j j j j �u����� ��u��"�M�� Qhp#j j j j �Q�������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rh#j j j j � �����(��u��-�M�QR�E�� P�M�Qh�"j j j j �ш���� ��u��E�    �G����E������   �j脜����ËE܋M�d�    Y_^[��]ÍI /���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    ���E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h�%j hy  h(j�Z�������u̃}� u0�s����    j hy  h(h�%h�%蒠�������sj�E������E�    ���M�}�t7�U��t��/   ��E��%��  ��/��/    �M���E������   �j������ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��j�h@�h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E��}� u!h�'j h�  h(j���������u̃}� u+������    j h�  h(h�'h�'�������s����u�fj�Å�����E�    ��/�E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j蛘����ËM�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��3��} ��]����������������̋�U��} u3��1j j �E�� P� �������u3���M�� Qj ��1R�,b]������������������������������̋�U��j�h`�h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP��������u3���   j�������E�    �M�� �M��U��B%��  ��t"�M��yt�U��B%��  ��t	�M��yukj�UR�EP���������tU�M��Q;UuJ�E��H;�<�} t�U�E��H�
�} t�U�E��H�
�} t�U�E��H�
�E�   ��E�    �E������   �j�Y�����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U��Q�EP蝃������u�����M�� �M��U��B��]������������������̋�U��Q��/�E��M��/�E���]������������������̋�U���/]����̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E܃}� u!h�(j h�  h(j蠀������u̃}� u.蹣���    j h�  h(h|(h�(�ؚ�����m  j荁�����E�    �U��/��E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡ�/�E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�Rh0(j j j j ������ ��u���M�Qh(j j j j �������u������E��/�H,�U��/�B0�E������   �j�^�����ËM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E�}� u!h�(j h�  h(j�"~������u̃}� u0�;����    j h�  h(h)h�(�Z�����3��  3҃} �U��}� u!h�(j h�  h(j�}������u̃}� u0�Ҡ���    j h�  h(h)h�(������3��0  3Ƀ} ���M�}� u!h�(j h�  h(j�P}������u̃}� u0�i����    j h�  h(h)h�(舗����3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u����t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M�谊���M��0{��P�MQ�#   ���M�蒟����]��������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E�    j�]|�����E�    h@*h� j j j j �{������u̃} t�M��U��/�E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u����u��  �U�z twj j�E�HQ��������tj�U�BP�0b��t$�M�QRh(*j j j j ��z������u��)�M�QR�E�HQh*j j j j �z������u̋E�HQh*j j j j �{z������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph�)j j j j �-z���� ��u̃=�/ t,j�U�� R�0b��u�E�HQ�U�� R��/����E�P�MQ�  ���   �U�zu;�E�HQ�U�� Rh�)j j j j �y������u̋M�Q�UR�x  ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Phd)j j j j �Uy���� ��u̋U�R�EP�  ��������E������   �j��������hH)h� j j j j �y������u̋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���t�h3ŉE��EP�M�荆���E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M���v����t3�M��v������   ~ �M��v��PhW  �E�P萓�����E��hW  �M�Q�M��v��P�Fr�����E��}� t	�U��U���E�    �E��M��L�������U��ڙ���     �E�Ph$�M�k��1   +�R�E�k��L�Q��������}*j h	  h(h�*hl*j"j膙���R�s���� �v����M��������U��D� �E�P�M�QhX*j j j j �v������u̍M������M�3��?�����]������������������������������������������������������������������������������������������������������������������̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP�4����E]������������������̋�U���8�h3ŉE��E�P�|�����}� u�}� u����t7�}� t1h�*h� j j j j �qu������u�j �(������   �3��M�3�������]������������������������������������̋�U���3��} ���E��}� u!h�(j h�	  h(j�jt������u̃}� u.胗���    j h�	  h(hH+h�(袎�����   �E�    �	�U����U��}�}>�E���<Q�U��E�L�Q�U��E�L�Qh$+j j j j �it���� ��u�볋E�H,Qh�*j j j j �Et������u̋E�H0Qh�*j j j j �#t������u̋�]�������������������������������������������������������������������̋�U��j j j �EP�MQ�$t����]�������������������̋�U��EP�MQj �UR�EP��s����]���������������̋�U��j j j �EP�MQ�UR�Rs����]���������������̋�U��j j j �EP�MQ�UR�EP�����]�����������̋�U��EP�MQj �UR�EP�MQ��r����]�����������̋�U��EP�MQj �UR�EP�MQ�UR�~����]�����������������������̋�U��j j �EP�MQ�UR��r����]�����������������̋�U���(�E��#E������E�u!h,j h�
  h(j�q������u̃}� u0�Д���    j h�
  h(h�+h,������3��@  �} t�U;Ur	�E�    ��E�   �E܉E��}� u!h|+j h�
  h(j�6q������u̃}� u0�O����    j h�
  h(h�+h|+�n�����3��   �}v�U�U���E�   �E؃��E3�+M���M�U�E�L�M��UU��U�E;E�v�ؓ���    3��i�MQ�URj�E�P�l�����E�}� u3��F�M�M�M�U��#�+M�M��E�+E���E�j��Q�U���R�G������E��M��E���]������������������������������������������������������������������������������������������������������������������������̋�U��j j �EP�MQ�UR�EP� p����]�������������̋�U��j j �EP�MQ�UR�EP�MQ��{����]���������̋�U���4�} u!�EP�MQ�UR�EP�MQ�%p�����  �} u�UR������3��  �E������E�j��Q�U��R�V�������t1�EPh�,j j j j�\o������u�������    3��C  j��R�E���P��������u�MQht,j j j j�o������u̋E��#E������E�u!h,j h�  h(j�Qn������u̃}� u0�j����    j h�  h(h0,h,艈����3��  �} t�U;Ur	�E�    ��E�   �EԉE؃}� u!h|+j h�  h(j��m������u̃}� u0�����    j h�  h(h0,h|+������3��  �U��P�O|�����M��U++E�}v�E�E���E�   �MЃ��M3�+U���U�E�M�T�U�EE�E�M;M�v�W����    3��   �UR�EPj�M�Q�}h�����E��}� u3��   �U�U�U�E��#�+U�U��M�+M���M�j��R�E���P��������M��U���E�;Ev�M�M���U�ŰE�P�MQ�U�R��z����j�E��Q詁�����E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es袎���    3��s�E�E�E��} t�MQ�UR�EP躇�����E��M Q�UR�EP�MQ�U�R�EP�k�����E�}� t �M�;M�s�U�+U�Rj �E�E�P��������E��]��������������������������������������������������������̋�U��EP討����]�������������̋�U��Q�} u�   �E������E�j��Q�U��R���������t!�EPh-j j j j��j������u��Lj��R�E���P��������u�MQht,j j j j�j������u�j�E��Q�$������]�����������������������������������������������������̋�U��Q���E��M���E���]������������������̋�U��Q��/�E��E���]�����������̋�U���/]����̋�U��EP�MQ�UR�h����]���������������������̋�U��� �E�    �E�    �E�    �E�    �E�    3��} ���E�}� u!h�-j h�  h(j��h������u̃}� u.������    j h�  h(hl-h�-����������w�E�    �U������U��E��Q�Ew�����E��U��E+�E�3�+M���M�}v�U�U���E�   �E����E�M�U�D
+E�E�M�+M�+M�M��E���]�������������������������������������������������������������������̋�U��Q�=  th �Ʉ������t�EP� ����z��h4�h��E������E��}� t�E��Gh$��,�����h�h ��R  ���=U thU�^�������tj jj �U3���]���������������������������������������������������̋�U��j j �EP�>  ��]���������̋�U��j j�EP�  ��]���������̋�U��jj j �   ��]�����������̋�U��jjj ��  ��]�����������̋�U���/����EP�Hj����h�   �i��]��������������̋�U��Q� 0�E��	�M����M��}� t�U��: tj�E��Q�T{������j� 0R�A{����� 0    �0�E��	�M����M��}� t�U��: tj�E��Q�{������j�0R��z�����0    j�0P��z����j�0Q��z����j�UR��aP�z�����0    �0    �n���U�8P�$b��u'�=8tj�8Q�ez�����8�8R�b��]�����������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    ��{���E�    �=80�U  �40   �E�00�} ��   �UQ��a�E�}� ��   �UR��a�E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�l���U�9u��E�;E�s�h�M؋R��a�E��gl���M؉�U܋UR��a�EСUP��a�E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���hL�h8��A  ��hT�hP��/  ���=<0 u#j��I������� t�<0   蹉���wv���E������   ��} t�6���Ã} t��80   �����MQ�f�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������̋�U���h�-�b�E��}� th�-�E�P��a�E��}� t�MQ�U���]�����������������̋�U��EP�������MQ�4b]�������������������̋�U��j��b����]���������������̋�U��j�v����]���������������̋�U��Q�(j���E��E�P�������M�Q老�����U�R�o�����E�P��[�����M�Q�d�����U�R�n������]����������������������̋�U��E;Es�M�9 t�U��ЋM���M��]�����������������������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�����������������̋�U���3��} ���E��}� u!h�.j h�  h@.j�Z`������u̃}� u0�s����    j h�  h@.h.h�.�z�����   �y3҃=,0 �U��}� u!h�-j h�  h@.j��_������u̃}� u0�����    j h�  h@.h.h�-�&z�����   ��M�,0�3���]������������������������������������������������������������������̋�U���3��} ���E��}� u!h�.j h�  h@.j�*_������u̃}� u0�C����    j h�  h@.h/h�.�by�����   �y3҃=(0 �U��}� u!h�.j h�  h@.j�^������u̃}� u0�ׁ���    j h�  h@.h/h�.��x�����   ��M�(0�3���]������������������������������������������������������������������̋�U���p�E�P�Hbh�   h /jj@j �������E��}� u�����  �M�� T��S    �	�U���@�U�� T   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M���S;U���   h�   h /jj@j ��~�����E��}� u��S�E��   �M��U��� T��S�� ��S�	�M���@�M��U��� T   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R�Db��t[�E����M������ T�M��U��E���
�U��E���Jh�  �U���R�@b��u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M��� T�M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P�<b�E��}����   �}� ��   �M�Q�Db�E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�@b��u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A�������SR�8b3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �	�E����E��}�@}y�M��<� T tg�U��� T�E��	�M���@�M��U��� T   9E�s�M��y t�U���R�Lb��j�E��� TQ�m�����U��� T    �x�����]���������������������������������������������������̋�U����=U u����E�    ��/�E��}� u����e  �M����t,�E����=t	�U����U��E�P��[�����M��T�U���juh00jj�E���P��y�����E�M�0�=0 u�����   ��/�U��	�E�E��E��M������   �E�P�[�������E��M����=��   j~h00jj�E�P�Py�����M��U�: uj�0P�Tl�����0    ����rj h�   h�/h�/h\/�M�Q�U�R�E�Q�{����P�g�����U���U��B���j��/P��k������/    �M��    � U   3���]��������������������������������������������������������������������������������������������������������������������̋�U����E�    �=U u�}���T1 h  hP0j �PbhP0�-~�����= U t� U���t� U�U���E�P0�E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   hl0j�M��U���P��P�����E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�   ���U����0�E��03���]�������������������������������������������������������������������������̋�U��E�(0]�����������������̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�h������t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P�>f������t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R��e������t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �Xb�E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j ��a�E��}� tjJh�0j�M�Q�IK�����E�}� u�U�R�Tb3��Dj j �E�P�M�Q�U�R�E�Pj j ��a��uj�M�Q�d�����E�    �U�R�Tb�E��]������������������������������������������������������������������������̋�V�����=(�s���t�Ѓ���(�r�^����������̋�V�0���=��s���t�Ѓ�����r�^����������̋�U��Q�E�   j h   j �\b��1�=�1 u3���   ��]�������������������������̋�U�졌1P�`b��1    ]�������������������̋�U��=�1 uhX1j jhh�0j�)N������u̡�1]�������������̋�U���0�E� �E�   �E���E��M����M�U��B3h�EԋM�Q�U�R��  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M���O���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=t� t ht��j������tj�UR�t����M����U�Hk���E��H;M�thh�U�R�M����U��<U���E��M�H�U�R�E�P��   ���U�M�I�s�������&�U��z�thh�E�P�M����������T���E��M߅�t�U�R�E�P�   ���E��]������������������������������������������������������������������������������������������������������������������������̋�U����E�8�t%�M��E��M��U�EB3E��E��M���r���M�Q�E��M��U�EB3E��E��M��r����]���������������������������������̋�U����E�    �E�    �=hN�@�t�h%  ��t�h�щl�   �U�R�pb�E��E�M�3M��M��lb3E�E���a3E�E��hb3E�E�U�R�db�E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M�h�U��҉l��]����������������������������������������������������������������̋�U��}csm�u�EP�MQ��g������3�]����������̋�U����qF���E��}� u3���  �E��H\Q�UR�S  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  � 2�U��	�E����E�� 229M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��;Ut�E����E��2k�M9M�s�ڋ2k�U9U�s
�E��;Mt3���E���]������������������������̋�U���(  ��2��2��2��2�5�2�=�2f��2f��2f��2f�|2f�%x2f�-t2���2�E ��2�E��2�E��2��������1  ��2��1��1	 ���1   �h�������l��������a��1j�O����j ��bh02�|b�=�1 u
j�iO����h	 ��xbP�tb��]����������������������������������������������������������������������������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh(3j jph�2j�iE������u̃}� u.�h���    j jph�2h�2h(3�_��������)  �} t�} u	�E�    ��E�   �M̉MЃ}� uh@2j jsh�2j��D������u̃}� u.�h���    j jsh�2h�2h@2�*_��������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�oW�����E��} u�E��P�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj ��^�����EċE���]�������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�b����]���������������̋�U��} u�T5    ��EP��a��S�T5   ]��������������̋�U���`�h3ŉE��E� �E� �E� �E� �E� �E� �E���E��E���E���E���E���E���E���E���E��E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E���E���E���E���E���E���E���E���E���E���E� �E� �E� �E� �E� �E� �E� �E׀�=T5 t��SP��a�E���E����M��M؋U�U��}��  4�}��  ��  �E����E��}��   ��  �M����M	�$�xM	�E�-�  �E��}���  �M��$�`N	�E�   �E� 4�U��]��E� �]��M��]ȍU�R�U؃���u�d��� "   �E�E���c  �E�   �E� 4�M��]��U��]��E� �]ȍM�Q�U؃���u�id��� !   �U�E���  �E�   �E�4�E� �]��M��]��U��]ȍE�P�U؃���u�d��� "   �M�E����  �E�   �E�4�U��]��E� �]��M��]ȍU�R�U؃���u��c��� !   �E�E���  �E�   �E�4�M��]��U��]��E� �]ȍM�Q�U؃���u�c��� "   �U�E���3  �E�   �E�4�E� �]��M��]��U��]ȍE�P�U؃��M�E����  �E�   �E�4�U�����  �E�   �E�4�E� �]��M��]��U��]ȍE�P�U؃���u��b��� "   �M�E���  �E�   �E�4�U��]��E� �]��M��]ȍU�R�U؃��E�E���S  �E�   �E�4�M��]��U��]��E� �]ȍM�Q�U؃���u�Yb��� "   �U�E���  �E�   �E�4�E� �]��M��]��U��]ȍE�P�U؃���u�b��� !   �M�E���  �E�   �E�4�U��]��E� �]��M�����U��E� �]��M��]��U��]ȍE�P�U؃���u�a��� !   �M�E���O  �E�   �E�4�U��]��E� �]��M��]ȍU�R�U؃���u�Ua��� !   �E�E���  �E�   �E� 4�M��]��U��]��E� �]ȍM�Q�U؃���u�	a��� !   �U�E���  �E�   �E��3�E� �]��M��]��U��]ȍE�P�U؃���u�`��� "   �M�E���k  �E�   �E� 4�U�����E��M��]��U��]��E� �]ȍM�Q�U؃���u�a`��� !   �U�E���  �E�   �E�4�E� ����M��U��]��E� �]��M��]ȍU�R�U؃���u�`��� !   �E�E���  �E�   �E�4�M�����U��E� �]��M��]��U��]ȍE�P�U؃���u�_��� !   �M�E���W  �E�   �E��3�U�����E��M��]��U��]��E� �]ȍM�Q�U؃���u�M_��� !   �U�E����  �E�   �E��3�E� ����M��U��]��E� �]��M��]ȍU�R�U؃���u��^��� !   �E�E���  �E�   �E��3�M�����U��E� �]��M��]��U��]ȍE�P�U؃���u�^��� !   �M�E���C  �E�   �E�4�U��]��E� �]��M��]ȍU�R�U؃���u�I^��� !   �E�E����  �E�   �E��3�M�����U��E� �]��M��]��U��]ȍE�P�U؃���u��]��� !   �M�E���  �E�   �E� 4�U��]��E� �]��M��]ȍU�R�U؃���u�]��� !   �E�E���O  �E�   �E�4�M��]��U��]��E� �]ȍM�Q�U؃���u�U]��� !   �U�E���  �E�   �E��3�E� �M�M��U��]��E� �]��M��]ȍU�R�U؃���u��\��� !   �E�E���   �E�   �E��3�M��M�U��E� �]��M��]��U��]ȍE�P�U؃���u�\��� !   �M�E���T�E�   �E��3�U��M�E��M��]��U��]��E� �]ȍM�Q�U؃���u�M\��� !   �U�E���M�3��E`����]ûD	E	SE	�E	�E	7F	�F	�F	tF	G	cG	�G	gH	H	�H	jM	 	
�I [I	�I	J	oJ	�J	'K	sK	�K	L	gL	�L	M	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E���#�S��S��S]������������������̋�U��j
��b��S3�]����������̋�U���h��  �,P��>�����E��M���  ���  ��   ���E�$�q9�����E�}� ~C�}�~�}�t�5h��  �U�R�>�����E��   �E�P���E�$j�^7�����   �M�Q�E������$���E�$jj�N3�����}���E�$�7�����]��E��E������Dzh��  �U�R�>�����E��D�B�E��� th��  �M�Q��=�����E��$�"�U�R���E��$���E�$jj��2������]������������������������������������������������������������������������������������̋�U��j
��b��S3�]�����������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������������������������������������������������������̋�U��=�  u0�EP���E�$�����$���E�$�MQj�vG����$�!��U��� !   h��  �UR�<�����E]���������������������������������̋�U����E�E�]��=�  u1�EP���E��$���E�$���E�$�MQj��F����$�!��T��� !   h��  �UR�;�����E���]����������������������������������̋�S�܃������U�k�l$���   �h3ŉE��C P�KQ�SR�S������u)�E�����E��KQ�SR�CP�KQ�S R�E�P�;�����KQ�xS������|����=�  u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q��E����$�%���|���R�7����h��  �C P�y:�����C�M�3��jW����]��[��������������������������������������������������������������������������̋�S�܃������U�k�l$���   �h3ŉE��C(P�K Q�SR�]R������u;�E����E��M������M��C�]��S R�CP�KQ�SR�C(P�M�Q�9�����SR�&R������|����=�  u?��|��� t6�C(P���C �$���C�$���C�$�KQ��|���R�D����$�%���|���P�I6����h��  �K(Q�&9�����C �M�3��V����]��[�����������������������������������������������������������������������̋�U����E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U�������������M�Q���ЋE�P�M�����҃������E�H���ʋU�J�E�����Ƀ������U�B�����M�A�U�������������M�Q���ЋE�P�M��� ��҃����E�H���ʋU�J�!;���E��E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E���t�M�Q���E�P�M��� t�U�B���M�A�U�%   �E�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�M����E��1�M�������E���M�������E���M�����E��M���   �U�t5�}�   t�}�   t�1�E����U�
�"�E������U�
��E������U�
�E%�  ���M��� ��ЋE��}  tT�M�Q ���E�P �M�Q ���E�P �M�U��Y�E�H`���U�J`�E�H`���U�J`�E�M��XP�X�U�B ���M�A �U�B �����M�A �U�E� �Z�M�Q`���E�P`�M�Q`�����E�P`�M�U��YP�/M���EPjj �M�Q��a�U�B����t�M�����E��M�Q����t�E�����U�
�E�H����t�U�����M��U�B���t�M����E��M�Q��t�E���ߋU�
�E����M�}�wb�U��$�]	�E���������   �U�
�@�E���������   �U�
�(�E���������   �U�
��E��������U�
�E������M�t�}�t�}�t.�;�U�%����   �M��%�U�%����   �M���U�%�����M��}  t�U�E�@P���M�U�BP���]�}\	e\	M\	5\	�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR�3����]�����������������������̋�U��j�EP�MQ�UR�EP�MQ�UR�e3����]�����������������������̋�U���D�E���E��M��t �U��tj�F;�����E�����E��  �M��t �U��tj�;�����E�����E��s  �M���   �U���  j��:�����E%   �E��}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z�H�]���H���]؋U�E���   �E�������z�H�]���X���]ЋM�E���Z�U�������z�X�]���H���]ȋE�E���,�M�������z�X�]���X���]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�%�����]�M��   �M��}�����}�E�����]��E�   �   ���]�����Au	�E�   ��E�    �U��U��E��f�E��M��f�M��	�U����U��}����}:�E��t�}� u�E�   �M���M�U��t�E�   ��E�M���M�봃}� t�E����]�U�E����E�   �}� t
j�8�����E�����E��M��t�U�� tj �8�����E����E�3��}� ����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �EP�  ���E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R�-�����E�P�bD������u�MQ�*�����E��"� h��  �U(R�o-�����EP�u*�����E ��]�������������������������������������������������̋�U��Q�E�E��}�t�}�~ �}�~���E��� !   ���E��� "   ��]��������������������̋�U��Q�E�    �	�E����E��}�}�M���0;Uu�E���4���3���]�������������������������������̋�U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]���������������������������������������̋�U����E�]��E�  �E��M���  �U����f�M��E���]��������������������������̋�U��Q�E%�  ��f�E��M����  f�M��E���]��������������������̋�U���E%�  ���ȋU�����P���E�$�+D����]��������������̋�U����E�]��E%�  �M���f�E��E���]����������������������̋�U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]�������������������������������������������̋�U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U�U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$�\B�����]��.j ���E�$�DB�����]��U���  ����-�  �E��M�U���E���]�������������������������������������������������������������������������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]������������������̋�U����E��t
�-x�]���M��t����-x�]������U��t
�-��]���E��t	�������؛�M�� t���]����]�������������������������̋�U��Q�=�S t�]���E�    �E���]�������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e�=�S ��   �E��@tp�=� tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe���    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]�������������������������������������������������������̋�U��Q�=�S t�]��e���U���]�����������������̋�U��Q�=�S t�����E��E���?�E���E�    �E���]����������������̋�U��Q�=�S t����E��E���?�E��(-����E�    �E���]���������������������������̋�U����=�S t8�>���E��E#E�M��#M���E��U������U��U��E�P�������E�    �E���]�������������������������̋�U��Q�����E��E��?E��E��M�Q�6������]�����������������������U���0���S�ٽ\�����=�  t�'-����8����   [����ݕz������U���U���0���S�ٽ\����=�  t��,����8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����,���   [�À�8�����=�/ uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��4������������4����s4��4�,ǅr���   ��4������������4����v��4VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P��%����_^�E�����U���0���S�u�u�   ���ٽ\�����8�����+������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[������������������������������������������������������������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^�����4�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����4�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����4���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�4��p��� ƅp���
��
�t������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    ����t
j
�-�����b���E��}� t
j�)��������tjh  @j�3����j�m����]��������������������������������̋�U��Q���E��M��#M��U#Uʉ��E���]���������������������̋�U��j�W,������tj�H,������u#�=�/uh�   �V����h�   �I����]�������������������������̋�U��Q�E�    �	�E����E��}�s�M��U;�(?u�E���,?���3���]�������������������������������̋�U���   �h3ŉE�EP��"�����E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j����������������� t������t���E�   ��E�   �}� ��  j�+������tj��*��������   �=�/��   j��<b�E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P������P������Q�U�R��b��  �}�   ��  ǅ�����5������-`5���  +ȉ�����������������j h  h8DhDhHChCh  h`5�6����P�m"����3�������f��  h  ������Rj ��b��u:j h  h8DhDhpBh8B������P������Q�36����P�"����������R�P��������<vk������P�9�����������TA�������j h  h8DhDh�Ajh�A������+�������������+�Q������R�G1����P�!����j h  h8DhDh Ah�@h  h`5��
����P�T!����j h  h8DhDhX@�E�Ph  h`5��
����P�!����h  h @h`5�8�����M�3��8����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �h3ŉE�}��  �E�E���p����M�ǅd���    ǅh����   ��h���R�E�P�MQ�UR�EP�������l�����l��� ��   � b��zt�  j j �MQ�UR�EP�]������h�����h��� u��   j^h�Ejj��h���Q�@1�����E��}� u��   ǅd���   ��h���R�E�P�MQ�UR�EP��
������l�����l��� u�   jih�Ejj��l���Q��0�����U���E��8 u�]j jlh`Eh4Eh�D��l�����Q�U�R��l���P�M��R������P�������d��� tj�E�P�#����3��-  ��d��� tj�M�Q�y#��������  �  �}��   �U��\�����\����     j j �MQ�UR��b��`�����`��� u�Zh�   h�Ejj��`���P��/������\������\����: u�(��`���P��\����R�EP�MQ��b��u�3��mj��\����P�"������\����    ����I�D�} u>ǅX���    j��X���R�E    P�MQ��b��u�����U��X����3������M�3��g4����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E��<]�����������������̋�U��E�U��DV�u�     j�E�P3�NVf�
��b��u3�^��]ËM�U�E�QRP��b��t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=�< u �=�< uH�  ��<��t:��<���<h\FP��a3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�RhXFV�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ��bP��b�����   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ��bP��b�M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �h3ŉE��=�< t3��M�3���/����]���<��   ����   VWh0F�b�= b�5�b��t?h  ������QP�օ�t,h  ������R������P��  ����t������Q�ׅ�uBh  ������Rj �օ�t,h  ������P������Q�  ����t������R�ׅ�u3�_^�M�3��-/����]����������������������������������������������������������������̋�U���  �h3ŉE�VhLG� b����u^�M�3��.����]�W�=�ah<GV�׉�������u_^�M�3��.����]�Sh(GV�׋؅�t4hGV�׋���t&������Pjj h�Fh  ���������tV��b[_3�^�M�3��8.����]Í�����Q������������R������Pj hpFQǅ����  �Ӌ�����R����V��b��u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M����F�F��E������F�H� F�P�$F�H�(F�Pf�,F�Hf�P������P� b�M�[_3�^�3-����]����������������������������������������������������������������������������������������������������������������������̋�U���  �h3ŉE��EV�uh   ������Qh   ������Rh   ������Qj�U�RP��.����$��t3�^�M�3��Y,����]�hxG������j	P�O)������u�hlG������jQ�5)������u�������R������P�E������Q�U�RPV� ���M������3�@^��+����]��������������������������������������������������������������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uhPIj jah�Hj��������u̃}� u.�'���    j jah�Hh�HhPI�8��������h  3҃} �U؃}� uhtHj jbh�Hj�������u̃}� u.�&���    j jbh�Hh�HhtH����������  j������E�    ��S�M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H��Sj�U�R�������43�uhHj jh�Hj�������u��E������%���    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;�StM�U�z t�E�H�U���M��E�H�J�U��    �E��S�H��S�E��M��S�h�   h�Gjj�S������E�}� u�E�������$���    �L�U��    �E��S�H�=�S t��S�E��M��A   �E�   �U�E�B�M��S�E������   �j������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�G �����E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR�1����]���������̋�U��P  �>����h3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �Pb��u8j h<  h�Hh�MhPMh4Mh  ������Q�$����P������������U��E�P�l������@v]�M�Q�[�����U��D��E�j hE  h�Hh�Mh(Lj��Q�U�������+й  +�Q�U�R������P�&�����} t'�EP��������@v�MQ�������U�DÉE���!�����������!���     �}uǅ�����K�
ǅ������U���t�M�������
ǅ������U���t�}uǅ�����K�
ǅ������M���tǅ�����K�
ǅ������} t�E�������
ǅ������} tǅ����xK�
ǅ������} t�M�������
ǅ������} tǅ����lK�
ǅ������}� t�U��������'�} t�E�������
ǅ������������������}� tǅ�����G�
ǅ������} tǅ����`K�
ǅ�����������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U���GPh�Jh�  h   ������Q�$ ����D�E�}� }*j h`  h�Hh�Mhl*j"j�����R�k����� ������������}� }8j he  h�Hh�Mh@JhJh   ������R�!����P�����h  h�I������P�U#����������������uj�|����j�o���������u�   �3��M�3��C#����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uhPIj jah�Hj��������u̃}� u.����    j jah�HhXNhPI����������h  3҃} �U؃}� uhtHj jbh�Hj�)�������u̃}� u.�B���    j jbh�HhXNhtH�d��������  j�������E�    ��S�M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H��Sj�U�R�h�����43�uhHj jh�Hj��������u��E������6���    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;�StM�U�z t�E�H�U���M��E�H�J�U��    �E��S�H��S�E��M��S�h�   h�Gjj��������E�}� u�E���������    �L�U��    �E��S�H�=�S t��S�E��M��A   �E�   �U�E�B�M��S�E������   �j�S����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR������]���������̋�U��X"  ������h3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj ��b��u8j h<  h�Hh�RhHRh8Bh  ������R�R����P�+�����������E��M�Q�i�������@v`�U�R�X������M��TA��U�j hE  h�Hh�Rh(Lj��P�M�������+����  +���P�M�Q�T����P������} t'�UR���������@v�EP��������M�TA��U��}��� �������p���     �}uǅ����0Q�
ǅ����,Q�M���t�E�������
ǅ����,Q�M���t�}uǅ����Q�
ǅ����,Q�E���tǅ�����@�
ǅ����,Q�} t�U�������
ǅ����,Q�} tǅ�����P�
ǅ����,Q�} t�E�������
ǅ����,Q�} tǅ�����P�
ǅ����,Q�}� t�M��������'�} t�U�������
ǅ����,Q�������������}� tǅ�����A�
ǅ����,Q�} tǅ�����P�
ǅ����,Q������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M��HNRh Ph�  h   ������P������D�E�}� }*j h`  h�Hh�Rhl*j"j�i���Q������� �Y����������}� }8j hc  h�Hh�RhHOh�Nh   ������P�<����P�����h  h�N������Q�����������������uj�����j�����������u�   �3��M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�B�����E��E�    �E���]�����������������̋�U����E�    �E�    �	�E����E��}�$}Z�M��<ʹuK�U�k����<�E��Ű�M����M�h�  �U��հP�@b��u�M��Ͱ    3��뗸   ��]��������������������������������������̋�U����E�    �	�E����E��}�$}O�M��<Ͱ t@�U��<մt3�E��Ű�M��U�R�Lbj�E�P�\�����M��Ͱ    ��E�    �	�U����U��}�$}3�E��<Ű t$�M��<ʹu�U��հ�E�M�Q�Lb뾋�]��������������������������������������������������̋�U��j�h@�h5�d�    P���SVW�h1E�3�P�E�d�    �E�   �=�1 u���j������h�   ��������E�<Ű t
�   �   h  h�Rjj�������E�}� u�0���    3��   j
� ������E�    �M�<Ͱ uDh�  �U�R�@b��u"j�E�P�����������    �E�    ��M�U�Ͱ�j�E�P������E������   �j
������ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��E�<Ű u�MQ���������u
j������U�հP��b]�����������������̋�U��E�ŰQ��b]��������̋�U��EPj ��bh�   ������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uhpTj jh�Sj��������u̃}� u0�0���    j jh�Sh�ShpT�R�����   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U�E�Ph�   �M��Q�}����3҃} �U��}� uh�Sj jh�Sj�R�������u̃}� u0�k���    j jh�Sh�Sh�S������   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U��E�Ph�   �M��Q�y�����tS��t3�t	�E�   ��E�    �M܉M�}� uh,Sj jh�Sj�7�������u̃}� u-�P��� "   j jh�Sh�Sh,S�r�����"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9�s
���E���M+M����U+щU؋E�Ph�   �M+M��U�D
P�����3���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��������������������������������������̋�U��j�h`�h5�d�    P�ĘSVW�h1E�3�P�E�d�    �} u3��   j���������u3��oj��������E�    �EP�MQ��>��	���URj �EP�MQ�UR�M�����M������E乀>� ����E������   �j�������ËE�M�d�    Y_^[��]��������������������������������������������������������������̋�U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� �����������������̋�U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]�������������������̋�U��j�h��h5�d�    P�ĘSVW�h1E�3�P�E�d�    �} u3��   j�
�������u3��pj�5������E�    �EP�MQ��>�&���U R�EP�MQ�UR�EP�M��E	���M��<
���E乀>�?����E������   �j������ËE�M�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�M��M������M���,�����E��>��>��>�} t�U��>�E��>���>    ��>    �M���,��>�U���>�E��>�M��>��> �E���]� ��������������������������������������������̋�U���H�M��M������M������=�> ��   ��>���?uG��>�B��@u8��>����>�U�R�6�����Ph]�E�P�q�����P�M�������v��>���?uS��>�H��$uEj �U�R������P�M������M������u��>��>�M�Q�������P�M�������U�R������P�M��w����M��p����u	3��  �?�M��Z����t������u��>���t��>R�M��M�����E�P�M��"����=�> u2�M���������>jh�>��>Q�������E��U���>�=�> ��   ��>P��>Q�M��������>�U�E�E�M����tY�E���� u0�U���U�E��  �M���M�U���� u�M���M�����U�E��
�U���U�E���E�띋M�U����>��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M�jPh�>�M�������>��]���������������̋�U���h�*�����tH��>%������>j �M�Q���������>��    ��>�E�P�M�����E�  �  ��>���?�t  ��>����>��>���?uK��>�H��?u=�U�R��������>���t��>����>��E�P�M�����E�9  �M�Q�������M������E�M��I����E��M��������u�U�R�M�R����E��  ��>�����   ��>���@��   �M�Q��	�����M���������   ��>��tn��> �E�P�M�Q�M����P�M��������>���@t>�M�Q�r	����P�M�������U�R�E�Ph$]�M�Q�M��A������l��P�M������)�U�R�E�Ph$]�M�Q�M��������A��P�M������}� t�M������}� t�M�������M�������u�M��w�����t�U�R�M�*����E��   �   ��>���t��>���@ut��>���t��>����>�5�����t:�}� u4�M�������u(�M��8���P�M�Q������U�R�M�����E�U��E�P�MQ�������E�>�j�M�����E�-�+��>���tj�M������E��j�M������E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�졠>���?uJ��>�B��$uj�MQ�R������E�;�$��>����>j j �EP�������E��j j�MQ�������E]�������������������������������̋�U���h�h3ŉE䡠>���0�M�x5�}�	/��>����>�E�P�MQ��>� ����E�;  �6  �M�� �����>���?ubj �M�Q�v�����P�M�������>���>����>��@t)��>����>��>�����ك�Q�M�����  jh@]��>R���  ����u�E�@]��>����>�9jh0]��>Q�ί  ����u�E�0]��>����>��E�    �}� ��   �E�P�������U�����twj�M�Q�M������U�R�(�����P��>���EЃ}� t�E�P�M������:h,]�M�����h(]�M�Q�U�R�E�P�M�Q��������������P�M��o����:h,]�M��K���h(]�U�R�E�P�M�Q�U�R������������P�M��3����N�E��t.��>���@u �M��7���P�M��������>����>�j@h�>�M������P�M������M��t��>�7�����u�U�R��>�1����E�P�M�c����E�M�3�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �M�������M�������E�    �E�    ��>��������>����>���������������_�o  ��������	�$�г	��>����>j�M�����E�  �M��u����M����   �U�R�p ����Pj<�E�P�	�����P�M��!����M������ȃ�>u
j �M��E ��j>�M��; ���} t�U���>���u�U�R�M�����E�  ��>����>��>�M�j j �U�R�������P�M��p����Eܣ�>�M�������u*��>�Q���1u�E�Pj~�M�Q�L�����P�M��2����M��{�����u�U�R�M��L����E�P�M������E�v  �%  ��>�Q����ZP�M������  �E�   ��>�Q����ZP�M��������  ��>��������>����>���������������_��  ���������	�$�L�	��>����>j�M������E��  ��>�B���@[Q�M��U����F  ��>�B���@[Q�M������E�  �  ��>�B���@[Q�M������M��p����U�R�M������E�F  ��  jh�Y�E�P��������M������M�Q�M�����E�  ��>�B���$[Q�M�<����E��  ��>�B���$[Q�M�����j j �U�R�������P�M��M����M�������u�M��r�����tj�M�����E�  �E�P�MQ�M������E�{  �  �  ��>�B���$[Q�M�������>���uj�MQ�M��o����E�4  ��>���0�E�x�}�rj�M�����E�  �M����\R�M�������>��������>����>�����������������0�����������>  ������$��	j �E�P�������M�Q�UR�E�P��t���Qj ��|���R�M��������� ����� ���E�^  �  �E�P�M�Q�M�� ��j,��d���R��l���P�������������P�M������j,��T���Q��\���R���������r���P�M�����j,��D���P��L���Q�y��������J���P�M�����j)��4���Rj ��<���P��������� ���P�M��i���j'�MQ�M��	����E�  �;�U�R�EP�M�������E�w  �!��>����>j�M�h����E�T  ��  ��>�B���$[Q�M��������  ��>��� �����>����>�� ��������������� t������0t!�N��>����>j�M������E��  j h\]�M�Q�������M��7����U�R�M� ����E�  j�M�����E�  �0  ��>���������>����>��������������������A������������	��   ����������	�$���	��>�Q����[P�M�^����E�  ��>�Q����[P�M��<�����>���?u5��,���P������P�M�������>���@u��>����>���$���Q�.�����P�M��_���hX]�M������U�R�M������E��j�M�����E�n�j�M�n����E�]�j�M�]����E�L�}� t
�M������-�M�������u!�E�PhxZ�����Q�!�����P�M������U�R�M�w����E��]ÍI �	2�	X�	~�	w�	��	n�	 �	�	&�	M�	��	��	��	ٮ	S�	X�	z�	<�	]�	 	

#�	p�	:�	:�	:�	��	��	        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�������>���>����>��@u��>���>����>��_tj�M�!����E�   ��>����>j �U�R�������j �E�P��������>���t��>���@t��>����>�ա�>���u��>����>j�M�����E���>����>�M�Q�M������E��]��������������������������������������������������������������������̋�U����   �M�������E� �M���������  ��>�����  ��>���@��  ��>��t��>��u�E�P�M�2����E�(  �M�������uE�M�Qh$]�U�R������P�M������E���t�M�Qj[�U�R������P�M�������E� ��>���?�  ��>����>��>���@�����@�����$��@�����@���%��  ��@�����T�	�$�@�	��>�B��_ua��>�Q��?uR��>����>�M�Q�U�Rj j �E�P��������������P�M��D�����>���@u��>����>�@�M�Q�U�Rj'�E�P�M�Q�9�����Pj`�U�R�������������������P�M��������   ��>����>�M�Q�U�Rj j�E�P�A��������h���P�M�������   j@h�>�M�������M�Qh\]�U�R�������P�M��{�����>�	�����u�E�P��>�����w��>����>�U�R��|���Pj]�M�Qj j�U�R�������������������P�M������E��*�E�P��l���Q��t���R�������������P�M�������.�E�P��\���Qj j��d���R�H��������o���P�M�����������>���<�����<��� t��<���@tW�W�M��������tj�M��?����;�U�R��D���Ph$]��L���Qj��T����������������������P�M��;�����
j�M�������U�R�M�����E��]Ðw�	��	¹	��	K�	 �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����>���uj�M�G����E�T�R��>���?u3��>����>j �U�R�������Pj-�EP�������E��j �MQ�������E��]�������������������������������������̋�U���   V�E�    ��>���Qu�E�x]��>����>��>���uj�M�y����E�S  �N  ��>���0��   ��>���9��   �}� tG��>� ��/��E��U���>����>�U�R�E�P�M�����P�M�Q�U�R��������E��4��>� ��/��E��U���>����>�U�R�E�P�M������E��M��M�U�R�M�����E�  �  �E�    �E�    ��>���@��   ��>���uj�M�r����E�L  �W��>���A|7��>���P*�E��U�������ȋ��>���A���M��u��j�M�����E��   ��>����>�e�����>���>����>��@tj�M������E�   �M��tX�}� t&�U�R�E�P�M�����P�M�Q�U�R�������E���E�P�M�Q�M��l����E��U��UЋE�P�M������E�V�T�}� t&�M�Q�U�R�M��N���P�E�P�M�Q�H������E���U�R�E�P�M��(����E��M��M��U�R�M�����E^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����>���u3���   ��   ��>���0|8��>���9*��>���/�M���>����>�E��   �   �E�    ��>���@tY��>���u3��k�7��>���A|$��>���P�U�����>��T
��U������2��>����>뚋�>���>����>��@t�����E���]����������������������������������������������������������������������̋�U����   ��>���?u��>�B��$tj�M������E�  ��>����>��>�U���>�E̋�>�M���\����#����M������M�������\�����>�E���>�MЉ�>�M��]����M��U����E� ��>���?u/��>����>�U�Rj��T���P�[�����P�M�������jj��L���Q�/�����P�M�袽���M��������t��>�U���up��D���P�������Pj<��<���Q�w�����P�M������M��y����Ѓ�>u
j �M�����j>�M������E��t��>���t��>����>�M���>�Ủ�>�E���>�M�Q�M������E��]�����������������������������������������������������������������������������������������������������������������̋�U���|�h3ŉE��E�   �M�������>�M��J������  ��>����  ��>���@��  �}� t	�E�    �
j,�M��v�����>���0�U�x4�}�	.��>����>�M�Q�U�R��>�0���P�M�������  ��>�E�M�������>���Xu��>����>h�]�M������%  ��>���$u7��>�H��$t)��>����>�E�P������P�M��D�����   ��>���?��   �E�P�)�����������tkj�M�Q�M������U�R������P��>���Eă}� t�E�P�M�������.h(]�M�Q�U�Rh�]�E�P�8��������8���P�M�诺���.h(]�M�Q�U�Rh�]�E�P������������P�M�������M������P�M�Q������P�M��_�����>+U��~��>�߼����u�E�P��>�ٹ���M�Q�M��Y����������> �U�R�M������E�M�3��b�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �h3ŉE衠>��M���>����>�E�������������R��  ��������$�	�$� �	�EP��������E�  ��>���@u$��>����>h�]�M�x����E�S  �3��D���Q�������P�URh����L����J������A����E�  �EP�������E�
  �M�Q�o������U�R�c������M����������   �M��������t{jd�E�P�M��6�����uj�M�����E�  �M��M��U���-u�E��E��E�.��E�.�M�Q�URje��4���P�M�Q��<���萸���������������E�]  �j�M�6����E�I  ��x���R�������=�����tSj��h���P��x���������h���Q������P��>����d�����d��� t��d���R�M�����E��  �E���Du5h(]�MQ��x���Rh�]��,���P�������������E�  �3h(]�MQ��x���Rhx]��$���P�^��������^����E�m  �h  j j ��\���Q�B����������R��������\���P�M�����E�/  j{��T���������M�������������H|3������J~�(�����R������P��T���腻��j,��T��������E���������������F������������wx�������$�x�	�����P������P��T����.���j,��T����_��������Q�������P��T�������j,��T����7���������R�������P��T����޺��j}�EP��T����{����E�-�+��>����>j�M������E�j�M������E�M�3�������]Ë���	Y�	m�	��	��	��	��	��	��	 �j�	B�	��	j�	B�	���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �M������
����E��M�����E��}���  uj�M������E�  �B�}���  u�EPj�MQ�������E�  ��}���  u�UR�M�����E�j  �E�% �  �0  �M��� �  t�U���   3���   ���������M��� `  ��Ƀ����������� t�U���   �� �����E�%   �� ����� ��� t>�M��� �  t�U���   3���   ���������
ǅ����    ������ ��
  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ t|�M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� @  tM�:�����t/�Է����t&�U�R�z�����Pj �E�P�Y�����P�M��?�����M�Q�T�����P�M��s����U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t�E�%   ��������M���   ������������ �-  �U��� �  t�E�%   3�=   ���������
ǅ����    ������ ��   �U�R�������P��|���Pj{�M�Q�M�:���������P�M��|����U�R�F������n�����u1h�^��l���P�M�Qj,��t���R�%�����������P�M��6���h�^�M������E�P������谳����tR�������tI�	�����u@�M�Q��T���Rj ��\���P�M�Qj ��d���R踿�������������K���P�M�萯���  �M��ٸ���M��Ѹ���M��ɸ���M�������M�蹸���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ �"  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t[�M���   ��   uJ��L���R������P�M�腮����D���P������P�M��m�����<���Q�}�����P�M��U����k�U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t'�E�%   =   u��4���Q������P�M�������,���R�������P�M��Э���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t8�U��� �  t�E�%   3�=   ���������
ǅ����   ������ u;�˴����t��$���R������P�M�����������P�������P�M�����蔰����tO�������t,�M�Q�����R�����P���������N���P�M�蓬��������Q������P�M�������������R�~�����P�M������M訿����uA�M�蜿����u)�w�����u �EPj ������Q�:�����P�M��R�����UR�M������E�    �M��Y����}� tNj ������P������Ph��������Q�P�����P�M�� ����������t�U�R�M�����E��  �bj h�>j������������������ t�������ڴ���������
ǅ����    �������E��M�Q������R�w�����P�M��M����E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ ��  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M���   ��   uzj,������R�E�P������Qj,������R�E�P������Qj,������R�E�Ph�^������Q���������������������������������������P�M��@����   �U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� tB�E�%   =   u3j,������Q�U�Rh�^������P���������n���P�M�跮���h�^�M�����h�^������Q�M�����P�M�苮��j)��x���R������P�#�����Pj(������Q�@�����������P�M��Q����U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� ��   �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t:�M��� �  t�U���   3���   ���������
ǅ����   ������ u�M�Q�M������̺����t��p���R�Q�����P�M��^������h���P�7�����P�M��]����]�����t�}� t�M�Q�M�������U�R�M������  �EP�M������M��� �  u.�U��� |  �� h  u�E�P�MQ�P������E��	  �1  �U��� �  u,�E�% |  = p  u�M�Q�UR芫�����E�	  ��  �E�% �  u]�M��� |  �� `  uLh�^�UR��X���P蠹����P��P���Qj{��`���R�M���������������萸���E�N	  �  �E�% �  u.�M��� |  �� |  u�U�R�EP�ڶ�����E�	  �[  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th�^�M������  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th\^�M��������   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tI�M��� �  t�U���   3���   ���������
ǅ����    ������ th ^�M��7����0�M��� �  u%�U��� |  �� x  u�E�P�M�\����E�  �M��� �  t�U���   3���   ����|�����M��� `  ��Ƀ���|�����|��� t�U���   ��x�����E�%   ��x�����x��� ��   �M��� �  t�U���   3���   ����t����
ǅt���    ��t��� u:�M��� �  t�U���   3���   ����p����
ǅp���    ��p��� t#�M�Qh����H���R������P�M��i�����E�P��@���Q迸����P�M��K����U��� �  t�E�%   3�=   ����l�����U��� `  ��҃���l�����l��� �x  ��������R  �E�% �  t�M���   3ҁ�   ��h�����E�% `  �������h�����h��� t[�M��� �  t�U���   3���   ����d����
ǅd���   ��d��� t!�M�Qh^��8���R�ٽ����P�M��W����E�% �  t�M���   ��   �s  �U��� �  t�E�%   3�=   ����`�����U��� `  ��҃���`�����`��� t�E�%   ��\�����M���   ��\�����\��� �$  �U��� �  t�E�%   3�=   ����X�����U��� `  ��҃���X�����X��� t�E�%   =   ��   �M��� �  t�U���   3���   ����T�����M��� `  ��Ƀ���T�����T��� t�U���   ��   tU�E�% �  t�M���   3ҁ�   ��P�����E�% `  �������P�����P��� t2�M���   ��   u!�U�Rh^��0���P�&�����P�M�褠���������  �M��� �  t�U���   3���   ����L�����M��� `  ��Ƀ���L�����L��� tl�U��� �  t�E�%�   3Ƀ�@����H�����U���   3���   ����H�����H��� t&�M�Qh�]��(���R�l�����P�M������Z  �E�% �  t�M���   3ҁ�   ��D�����E�% `  �������D�����D��� tp�M��� �  t�U����   3����   ����@�����M���   3ҁ�   ��@�����@��� t&�E�Ph�]�� ���Q踺����P�M��6����   �U��� �  t�E�%   3�=   ����<�����U��� `  ��҃���<�����<��� tb�E�% �  t�M����   ��Ƀ���8�����U���   ��҃���8�����8��� t!�E�Ph�]�����Q������P�M�苞���U��� �  t�E�%   3�=   ����4�����U��� `  ��҃���4�����4��� t�E�%   ��0�����M���   ��0�����0��� t*�O�����u!�U�Rh�]�����P�w�����P�M�������M���   t!�U�Rh�]�����P�K�����P�M��ɝ���M�Q�M衴���E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���x�E�    ��>���_u�U��� @  �U���>����>��>���A�  ��>���Z�  ��>���A�E���>����>�U��� �  �U��E���t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M�U����U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U��E��E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E܋M܉M��;�U��� �  t�E�%?����E���M��������M؋U؉U���E���  �E��k  �E����Eԃ}���   �M��$�8�	�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M̋ỦUЋEЉE����E���  �E��  �  ��>���$��  �E� ��>����>��>��Uȃ}�R�]  �E���|�	�$�T�	�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  ��>�Q��Pu��>����>��>����>��>��Eă}�Q��   �M�����	�$���	��>����>�1����  ��>����>��>���0|C��>���95��>���>�D
ѣ�>�����E��M���   �M��E��-  ��E���  �7��>����>读���	  �E���  �E���  �E���  �E���  ��  �E���  ��>����>��  �E���>����>��>���0|��>���5~$��>���t	�E���  ��E���  �E��z  ��>���0�E��M��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��M���t�U���    �U���E�%�����E��M����M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  ��>����>��  ��>���0��  ��>���8��  ��>��U졠>����>�M�������M��U�U��E���0�E��}��?  �M��$�8�	�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C��>���9u��>����>�E���  ���>���t	�E���  ��E���  �E���]ÍI n�	p�	�	p�	��	p�	��	K�	=�	��	��	��	(�	��	�	d�	�	 																																																																					�(�	��	��	�	7�	 ����	@�	��	i�	��	}�	��	��	��	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j ������P�M�������>���tl��>��E��>����>�U�U�}�0t�}�2t�}�5t(�5h�]�M�蕪���&�E�P������P�M������j�M�Y����E�(�
j�M�蜍��h�^�M��T����M�Q�M藡���E��]���������������������������������������������������̋�U���@�M�迓��j j�E�P�ݟ����P�M��P����M��I�����uN��>���tA��>���@t4�U�R�E�Ph$]�M�Q�U�R蜷������膛����豹��P�M��������>���@u��>����>�b��>���tj�M�艸���J�M��	�����tj�M��q����2�U�R�E�Ph$]�M�Qj�M��	������������1���P�M��v����U�R�M�N����E��]��������������������������������������������������������������������������̋�U�����>����  ��>���A�E���>����>�}���   j�M��K���蔌������   �U�����U��}���   �E�����	�$���	j�\�����P�M�記���|j�G�����P�M�蓘���gj�2�����P�M��~����Rj������P�M��i����=j������P�M��T����(j������P�M��?����j�ސ����P�M��*����U�R�M�����E� �j�M�l����E��j�M�[����E��]ÍI ��	��	��	��	�	$�	9�	L�	 ��������������������������������������������������������������������������������������������̋�U�졠>���@u"��>����>�EP�M�~����E���MQ�UR腇�����E]�����������������������̋�U��� �EP�M��7�����>��U��}� t�}�?tq�}�Xt��   �E�Pj�MQ�p������E��   ��>����>�M��ә����th�]�M�%����E�   ��E�Ph�^�MQ�ˡ�����E�w��>����>�E��j �M�胏��P�E�P�M�Q�U�R������P�M������E�P�MQ�������E�$�U�R�M�Ҝ���E��E�P�MQ�������E��]�������������������������������������������������������������������������̋�U���<�M��ώ����>��Mȃ}�B��  �U�����	�$���	�MQj�UR�������E�j  h_�M��I����M�u�����u
j �M�膰���EP�M�������>����>�E����U�R�M�这��P�E�P�MQ�������E�   ��>�B��$t<��>�Q��u�EPj�MQ�o������E��  �j�M�����E�  ��>����>��>��Mă}�T�o  �U����	�$���	��>����>�UR�EP菪�����E�Y  ��>����>j�UR�EP輆�����E�0  ��>����>�E�j �M��5���P�U�R�EP�M�Q藯����P�UR��������E��   ��   h_�M�������M������u
j �M�������EP�M��e�����>����>�E�4Z�U�R�M��6���P�E�P�MQ苲�����E�z��>����>j�M謝���E�\�G��>����>h_�M�Ã���E�;�&�MQj�UR�Ř�����E�"j�M�c����E��EP�MQ�������E��]Ë��	��	C�	 �	w�	 �Q�	
�	1�	Z�	��	��	�	0�	h�	 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� ��>��M�}�XtD�}�Zt�`��>����>������t	�E�G��E�<_�E�P�M�i����E��   ��>����>h�]�M�E����E��   �U�R�������M��v�������   ��>��M�}� t�}�@t`�}�Zt�v�U�R�M�'����E�   ��>����>�E�����t	�E�4_��E�$_�M�Q�U�R�M�腑��P�M������E�>��>����>�M�Q�M����E� j�M�K����E���U�R�M蠖���E��]��������������������������������������������������������������������������������������������̋�U���,�E�   �M�蘈���M��;������  ��>���@��   ��>���Z��   �}� t	�E�    �
j,�M��f�����>�����   ��>���0�M�x3�}�	-��>����>�E�P�M�Q��>����P�M��փ���k��>�U�M�����P�E�P螭������>+M��~��>������u�U�R��>��}���E�P�M��~�����>;M�u
j�M�������j�M�������������U�R�M������E��]����������������������������������������������������������������������������������������̋�U���(��>���tg��>���Zu'��>����>�M��ֆ��P�M�[����E�^�0j)�UR�E�P�@�����PhL_�M�Q�Ř�������%����E�,�*j)�URj�E�PhL_�M���}�����������������E��]�������������������������������������������������������̋�U���x��>����k  ��>��E���>����>�E� �E������M������U��U��E���C�E��}��   �M���H	
�$�	
h`�M��y����?  h`�M��g����-  h`�M��U����  h`�M��C����	  h `�M��1�����  h�_�M�����h�_�M�芛����  �E����E���  ��>��U��E�E���>����>�U��U��}�Y�8  �E����	
�$�h	
�E������(  h�_�M�裋���  h�_�M�葋���  h�_�M�������   h�_�M��m�����   h�_�M��[�����   h�_�M��I����   h�_�M��7����   h�_�M��%����   ��>����>�E�P�,�����P�M���z���M��(�����t�M�Q�M諑���E�~  �R�UR�E�P������Ph�_�MQ�������E�R  ��>����>j�M��A����h�_�M�舊���Qh�]�M��y����B��>����>�M�Q腄����P�M��8z���M�聍����t�U�R�M�����E��  �}����   �E��E��M���C�M��}���   �U���

�$��	
�M�Qhx_�U�R�G�����P�M���y���e�E�Phl_�M�Q�'�����P�M��y���E�U�U��E���E�E��}�w/�M���0

�$�(

�E�Phx_�M�Q�������P�M��^y���M觌����u�URj �E�P�Q�����P�M��i~���M�Q�M�����E��   ��   �M��l����UR�M������}��uF�M��:����E�P�M�Q�U�R�,������M��R�����uh�Z�M��d����E�P�M觏���E�}�M������tA�M���t$hd_�M�躈���U���thX_�M�������E���th_�M�莈���M�Q�U�R�EP�G������E���MQj�UR�������E��]��


&
8
W
J
i
�
x
�
   










	�I �
�
�
�
�

 
�
�
2
D
V
�
 	
���
v
�
�
 �I �
�
     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�;�����t�ȕ����u	�E�   ��E�    �EЉE��M���~����>��U̡�>����>�M̉Mȃ}�Y��   �U���$
�$�
��>����>he`�M��u���E�   h\`�M��#����khP`�M������\hH`�M������Mh<`�M�������>h,`�M������/�b����E��U�R�b�����Ph$`�E�P������P�M��t���M���}���}� t�M�Q�M��t���U�R�
w����P�M��y���E�P�M�B����E��]Ë�"
F
U
d
�
s
�
�
 ���������������������������������������������������������������������������������������������������������������������������������̋�U��EP�;������E]����������̋�U����M��|����>�����   ��>��E�M��0�M�}�wH�U��$�4
h�`�M������>h�`�M�������/�-hx`�M������h�_�M��Ղ���j�M�(����E�~��>��M��>����>�E�E�M��1�M�}�w/�U���\
�$�T
�M�Qhx_�U�R�ˍ����P�M��Ir���E�P�M�!����E��j�M訌���E��]�e
e
t
t
�
�
�
�
�

    ��������������������������������������������������������������������������������������������̋�U����   ��>���u�URj�EP�?������E�  ��>���6|��>���9~ ��>���_tj�M豋���E��  ��>���6�U���>����>�}�)u[��>���t2��>���=�M���>����>�}�|�}�~�E�������EPj�MQ艆�����E�M  ��}� |�}�~�E������}��uj�M�	����E�   �M���y���UR�M��U����E����  �M�Qh$]�U�R�ɋ����P�M��Gp����>���t5�U�R�E�P�M�Q趝����Pj �U�R�)��������ß��P�M��p����E�Pj�M�Q�Å����P�M���o����>���t1��>���@u��>����>�j�M�3����E�J  ��M�Qj�UR�j������E�.  �Tw����t�E�P藆����P�M��uo����M�Q耆����P�M�詒���U���tS�s����t5�E�P�M�Q�U�R�\|����Pj �E�P�;�������՞��P�M��o����M�Q�/|����P�M��N�����r����t)�U�R��x���P�M�Q���������莞��P�M���n�����p���R�؜����P�M������M������u.j)��`���P�M�Qj(��h���R�~�������h���P�M��n��j h�>j苆������\�����\��� t��\����w����0����
ǅ0���    ��0����E��M�Q�U�R�Jx����j)��D���P��T���Q������Pj(��L���R�~�������؜��P�M��!s���u����t�E���t�M�Q�M��s���Q�����t��<���R��|����P�M���r�����4���P�|����P�M������}� t�M�Q�M��m���j�M������E��U�R�M�L����E��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����>�����   ��>���6|��>���9~��>���_un�UR�M��l���M�E����u$�M�9����u�M�$�����u�EP�M���p���M�����u�MQ�M���p���U�R�EP�������E�   �>j �MQ�UR�EP�M�Q�M������U�3Ƀ�*��Q�U�R�EP�n�����E�m�kj�M��̅���MQ�M��ي���M�~����u�UR�M��^p���M�u~����u"�M�i~����u
j �M��z����EP�M��0p���M�Q�M�ց���E��]��������������������������������������������������������������������������������������������������̋�U���4�M���s����>����>��>��UЀ}�At�}�BtN�}�C��   �   �} u%�E����&u	�E����E�<Z�E�M̉��>����>�  �} tj�M�s����E�}  �E� j>�M��Ӊ����>����>�N  �U����>����>�3  ��>���t��>�H��uj�M�����E�  �} tj�M������E��   ��>���0����>�Q�DЉE��>����>�}�v/j,�M��!����U�3�PR�M�茇��P�M�Q�M��Ø��P�M��i��j>�U�R�M��ڗ��P�M���h����>���$u��>����>�j^�E�P�M�襗��P�M��h����>���t��>����>�
j�M��fk���M������M�Q�M�f���E��M��q���E��]�����������������������������������������������������������������������������������������������������������������������������������������������������̋�U���$  �M��q���E� ��>����  ��>���$u8�MQ�U�R�EP�M�Q�s�����M���z����u�U�R�M�X~���E�  ��>���>�3҃�A����+��+ʉM�M��p���M��p���E�   �E艅����������t������tw��������   �  ��j����tW踃����tN�M��8z����u/j�o����P�M�Qj �U�R�M�覕�����?x��P�M��f���j�ro����P�M��v���   �aj����tN�M���y����u/j
�Eo����P�E�Pj �M�Q�M��J�������w��P�M��Zf���j
�o����P�M��bv���`�j����tN�M��y����u/j	��n����P�U�Rj �E�P�M��������w��P�M��f���j	�n����P�M��	v����E�    �}� t|��>����>��>���$u8�MQ�U�R�EP�M�Q��q�����M���x����u�U�R�M�t|���E�  ��>���>�3҃�A����+��+ʉM�}� �)�����>���t��>����>�}���  �EP�M���e���M�Q�U�R�M��Ȕ��P�M��e���M��Vx����u)�E�P��|���Qj �U�R�M��ȓ����蓔��P�M���d���M��!x����u,�E�P��l���Qj ��t���R�M�萓�����[���P�M��d���E���  �} tj�M� ���E�  �M���tz�E�Ph$]��d���Q������P�M��Qd����>���t,�M�Q��T���R��\���P蹑�������Փ��P�M��d����M�Qj��L���R��y����P�M���c���$��>���t��D���R�l�����P�M�������>���uj�M��f���/��>���>����>��@tj�M�~���E�  �Rg����t[�U��������������t�B�} tj�M��}���E�t  �E�P��4���Q��<���R�^p����������P�M��+c���#�E����u��,���Q�2p����P�M��Q����U��t!�E�Ph�`��$���Q�_~����P�M���b���U��t!�E�Ph�`�����Q�6~����P�M��b���} ��   �M��u������   �M��y����u�M��u����t:�M��w����t�UR�M��jb����EPj �����Q�dr����P�M��|g���@�UR������Pj �����Q�URj �����P�0r��������������Ñ��P�M��:g���*�M�Ou����u�MQj ������R��q����P�M��g���M��v���E���t�M��6r���M�Q�M�x���E��   �j�M� |���E�   �   �} ux�M��t����ul�M��x����u�M��t����t�URj�EP�*w�����E�u�9�MQ�URj ������P�MQj������R��v�������������Ґ���E�:�8�} u%�M�\t����u�EPj�MQ��v�����E��j�M�`{���E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����>����  �} t]��>���XuO��>����>�M�'r����th�]�M�y_���E��   ��URh�^�EP�z�����E��   ��>���Yu%��>����>�MQ�UR�h�����E�   �EP�M�Q�x�����M�<a����t �U�Rh�`�E�P�y����P�M��1^���*�M�<v����t�M�Qh�`�U�R�y����P�M��^���E�P�M��t���E���MQj�UR�s�����E��]��������������������������������������������������������������������������������̋�U���   ��>����s  �l���E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M��z�����ه��������P�MQ�[w�����E�  �  �M��cf���M�wr����th�Z�M��|���M��ko����tR�U��E����E���tB��>���t5j]�E�Pj �M�Q��t����Pj[�U�R�l������聋��P�M���a��뢋M��o����u^�M��q����t�E�P�M�Q�M� ���P�M��e\���7�U�R�E�Pj)�M�Q�URj(�E�P�Tl����������������P�M��,\���M�Q�U�R�6������M��R����E�P�M��r���E�   �   �M�Do����uSj]��|���Qj�U�Rh�`�E�P�MQj(�U�R��k�������>m�����Z�����萊��P�EP��u�����E�?�=j]��d���Qj��l���Rj[��t�����x�����������O���P�EP�u�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j'�EPj �M�Q��r����Pj`�U�R�j�������w����E��]�����������������������̋�U����E��j�M��c��P�E�P�M��c��P�MQ�������E��]����������������������̋�U��Q�E�pZ�E�P�MQ�UR�EP�p�����E��]��������������������̋�U��Q�E���E�P�MQ�UR�EP�Vp�����E��]��������������������̋�U��EP�MQ�UR�EP�p�����E]��������������̋�U��j�EP�q�����E]��������̋�U��j �EP�q�����E]��������̋�U��j �EP�kq�����E]��������̋�U��EP�MQ�s�����E]������̋�U��Q��>��M��}� t)�}�At�0��>����>h�`�M�sY���E�j�M�,s���E�j�M�s���E��]���������������������������������̋�U���@�EP�M��Io���M���j�����b  ��>����Q  �E�P�M�Qj �U�R�E�P�:n�������������·��P�M��X���M��j�����  ��>���@��   h�`�M��yw���M��[j������   ��>�����   ��>���@txj'�M�Q�U�R�3�����Pj`�E�P�g�������n���P�M��\����>���@u��>����>�M���i����t��>���@th�`�M���v���Z����M��i����t ��>���u
j�M���Y��j}�M�肂����>���@u��>����>�'�M��ji����t�U�Rj�E�P�l����P�M���V���M�Q�M�m���E��]����������������������������������������������������������������������������������������������������������������̋�U��EP�W�����E]����������̋�U����E��j �M��f_��P�E�P�M��Y_��P�MQ�Á�����E��]����������������������̋�U����EP�M��l��h�`�M��Mu���M�Q�;�����P�M���Z��j}�M��	�����>���@u��>����>�U�R�M�Tl���E��]��������������������������������̋�U���,j h�>j�Mm�����E��}� t�M��u^���E���E�    �EԉE�M�Q�U�R�}U�����EP�M�Qj �U�R�E�P��j������較����臄��P�M���T���M�Q�M�k���E��]������������������������������������������������̋�U�조>�������]����������̋�U�조>%   �����]��������̋�U�조>�������]����������̋�U�조>�������]����������̋�U�조>�������]����������̋�U�조>��`3Ƀ�`����]�������̋�U�조>%�   �����]��������̋�U�조>%   �����]��������̋�U�조>%   �����]��������̋�U�조>%   ]���������������̋�U�조>%    ]���������������̋�U�조>% @  ]���������������̋�U�조>% �  �����]��������̋�U�조>%   �����]��������̋�U���X����t�E��H[���M��H[��]���������������������̋�U�조>�������]����������̋�U��EP�MQ��>�r��]�������̋�U����M�E������E�} t�MQ�U��Ѓ���   ��   �} w�E   �M�Q;U��   �}   v3��   jh�>h  ��i�����E��}� t�M��u���E���E�    �E��E��}� tA�M�y t�U�B�M���U�E��B��M�U��Q�E�M��H�   +U�E�P�3��!��M�Q+U�E�P�M�Q�E�H�D
��]� ���������������������������������������������������������������������̋�U��Q�M��E��     �E���]�������̋�U����EP�MQ�UR�M��+n�����g����E��]���������������������̋�U����EP�MQ�UR�M���j�����(����E��]����������������������̋�U����EP�MQ�UR�M���P���������E��]����������������������̋�U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]�����������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��f���E���]� ������������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��} tdj h�>j��e�����E��}� t�EP�M���S���E���E�    �M��U��E����Ƀ�������   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ���������������������������������������������������������������������������������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ��"  ���E��}� v�U�R�EP�M��9c���E���]� ���������������������������������������������������������������������̋�U���V�M�E�H�� ����U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E��     �M�Q�������E�P�M�Q�������E�P�M�Q�������E�P�M�Q������E�P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	�H����t�U����U���E�H�� ������U�J�   ������E�P�M�Q�M���`���U����t<�U�E���M�	���u�;�t�U�B% ������M�A�U��    �!�M���y����u�E�H�� ������U�J��E�H�� ������U�J��E�H�� ������U�J�E�^��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�조>%   ]���������������̋�U���$�h3ŉE��M܍E��E��M܋Q�� ����E܉P�M��    �U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%����M܉A�U�� �E����E�j j
�MQ�UR�po����0�� �M��j j
�UR�EP�Qm���E�U�MMu��U��E�+й   +�Q�U�R�M��6^���E܋M�3���r����]� ����������������������������������������������������������������������������������������̋�U���(�h3ŉE��M؍E��E܋M؋Q�� ����E؉P�M��    �U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%����M؉A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U܃��U�j j
�EP�MQ�m����0�� �U܈j j
�EP�MQ�k���E�U�UUu��E��t�M܃��M܋U��-�E܍M�+��   +�R�E�P�M��f\���E؋M�3��q����]� ��������������������������������������������������������������������������������������������������������̋�U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�h�����M���U��: u�E��H�� ������U��J�E���]� �����������������������������������������������������������������������̋�U��Q�M��E��H����3�������]���������������̋�U��Q�M��E�3Ƀ8 ������]������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J�E���]��������������̋�U��Q�M��E��@������]�������̋�U����M��M��WU����u�E��H��	��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��M��	U����u�E��H��   �U��J��]���������������������̋�U����M��M���T����u�E��H��
��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��    �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� @  �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� �  �U��J��]�����������������̋�U��Q�M��M���R����t3���E���U����ȋ�Ћ�]�����������������̋�U��Q�M��M��R����t2���E���U����ȋB�Ћ�]����������������̋�U����M�M��gR����uX�} u*�M���e�����Ej h�>�EP�W�����E��M��M�} t �U�E�L�Q�UR�M��P^���E��E��  ��} t�M� �E��]� �������������������������������������������̋�U��Q�M��M��Q����t�E��EP�MQ�U���M��	��B�Ћ�]� ����������������������̋�U����M�E�P�M���T���MQ�M��ui���U�R�M��T���E��]� ����������������������̋�U����M�E�P�M��T���MQ�M��K]���U�R�M�T���E��]� �����������������������̋�U����M�E�P�M��VT���MQ�M��B���U�R�M�>T���E��]� �����������������������̋�U����M�E�P�M��T���MQ�M��d���U�R�M��S���E��]� �����������������������̋�U����M�E�P�M��S���MQ�M��?���U�R�M�S���E��]� �����������������������̋�U����M��} t_j h�>j�T�����E��}� t�EP�M��R�M���Q���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ������������������������������������̋�U����M��M��UN����tb�E��tZ�M��O����t�MQ�M��[���?j h�>j�S�����E��}� t�UR�M���[���E���E�    �E�P�M��X���E���]� ���������������������������������������������̋�U����M��M��M����tu�} to�E���te�M��[N����t�UR�M��K���Kj h�>j�S�����E��}� t�EP�  ��P�MQ�M��K���E���E�    �U�R�M���W���E���]� ������������������������������������������̋�U��Q�M��M���L����tG�M�M����t�M�Qk��P�M��=���(�M��M����t�EP�M��-:����M�R�M��FW���E���]� ��������������������������̋�U����M��M��eL������   �} ��   �M��M����t�EP�M���B���j�M�j����t�M�j����u@j h�>j�Q�����E��}� t�MQ�M��?���E���E�    �U�R�M��V����M�Zj��P�M�� <���E���]� ���������������������������������������������̋�U��Q�M��M��K����tC�M��ML����u�}t�}u�EP�M��g����} u��MQ�^����P�M���U���E���]� ������������������������������̋�U����M��M��i����t3�M��J����u'�M�ni���E��E�%�   �M��Q�� ���ЋE��P�E���]� ���������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��O���E���]� ������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�  ��P�UR�M���M���E���]� ���������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h�>j�)M�����E��}� t�MQ�M��;���E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������̋�U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ��X�����U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ������������������������������������������������������������������̋�U����M�E�8 tj�M���a���  �} ��   �} ��   �M�M��}� t�}�t�u�U�B% ������M�A�   j h�>j��J�����E��}� t�U�P�M���R���E���E�    �M�U��E�8 u�M�Q�� ������E�P�[j h�>j�fJ�����E��}� t�MQ�UR�M���B���E���E�    �E�M��U�: u�E�H�� ������U�J��E�H�� ������U�J��]� ����������������������������������������������������������������������������������������̋�U��Q�M��E�3Ƀ8	������]������̋�U��Q�M��E�� �����E���]�������̋�U����M�M���3����uf�M�{D����uZj h�>j�2I�����E��}� t�EP�M���G���E���E�    �M��M��}� t�U����M��U��M�U��T��E��]� �����������������������������������������̋�U��Q�M��} |�}	~j�M��J���E�;�9�E��8�t
�M��U;~j�M��J���E���E�M��T�R�M�!G���E��]� ��������������������������̋�U��Q�M��E�� �`�E���]�������̋�U��Q�M��M���Q���E�� �`�M��U�Q�E���]� �������������������̋�U��Q�M��   ��]��������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E;Es�M�U��B��M���M�E��]� �����������������̋�U����M��M��Q���E�� �`�} tP�} tJj h�>�MQ�G�����E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ�S  ����U��B    �E��@    �E���]� ������������������������������������������������̋�U��Q�M��E��@��]�������������̋�U����M��E��x t�M��Q�E��H�T
��U���E� �E���]����������������������������̋�U��Q�M��E��HQ�U��BP�MQ�UR�/W������]� ������������������̋�U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�"  ���EE��]���������������������̋�U����M��M��XO���E�� a�} t#�M�P^����t�M�C^����u	�E�    ��M�M��U��E��B�E���]� ����������������������������������̋�U����M��E��x t�M��I��S���E���E�    �E���]��������������̋�U����M��E��x t�M��I�N���E���E� �E���]�����������������̋�U����M��E��x t�MQ�UR�E��H��K���E���M�M��E���]� ��������������������̋�U��Q�M��M��
N���E�� a�M��U�Q�E��H����Ƀ�����U��J�E���]� ��������������������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E��x��,"/a��]�����������������̋�U��Q�M��E��xujh,a�MQ�UR�T������E��]� ���������������������������̋�U��j�h�d�    P�h3�P�E�d�    �d?��uM�d?���d?�E�    j �(?�;Z��j�4?�/Z��j�@?�#Z��j�L?�Z���E������} |�}}�Ek�(?��L?�M�d�    Y��]��������������������������������������������������������̋�U��Q�M��M��*L���E�� 4a�M��U�Q�E��M�H�U��B�����E���]� ����������������̋�U��QV�M��E��x }.�M��Q�E��H���Ћ��M��Q�E��H������M��q�U��B^��]��������������������̋�U����M��E��H�U��B��ȋB�ЈE��M���u�U��B�M��I��B�ЈE��E���]������������������������̋�U����M��EP�MQ�U��B�M��I��B�ЉE��M�;Ms�UR�E�P�M��Q�E��H��B�����E���]� ����������������������̋�U��Q�E�    �	�E���E�M���t�E����E���E���]����������������������������̋�U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]��������������������������̋�U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]������������������������̋�U��Q�E�    �}�wC�EP�S�����E��}� t�*�=X5 u��O���    ��MQ��?������u����UR��?�����O���    3���}� u�O���    �E���]���������������������������������������̋�U��Q�=�1 u��G��j��/����h�   �/�����} t�E�E���E�   �M�Qj ��1R��b��]�������������������������̋�U��QV�E�    �} u�4�EPj ��1Q��b�E��}� u� bP�7�������N���0^��]���������������������������������̋�U��E�h?]�����������������̋�U��Q�h?�E��M�Q��a�E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�D����]����������������������̋�U��jh �j�I����h ��xbP�tb]����������������������̋�U���8  �h3ŉE��}�t�EP�3����ǅ����    jLj ������Q�<V�����������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M��������a�E�j ��b�U�R�|b���������� u�}� u�}�t�EP�2�����M�3��nP����]�������������������������������������������������������������������������������������������������̋�U��Q�E�    �h?�E��M�Q��a�E��UR��a�E�E�h?�E���]������������������̋�U��Q�E�    �h?�E��M�Q��a�E��E���]�����������������������̋�U��EP�MQ�UR�EP�MQ�B����]�������������̋�U��EP�MQ�UR�EP�MQ��A��]�����������������SVW�T$�D$�L$URPQQh0_
d�5    �h3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�A���   �C�_)���d�    ��_^[ËL$�A   �   t3�D$�H3��iN��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�A��3�3�3�3�3���U��SVWj Rh�_
Q�c7��_^[]�U�l$RQ�t$������]� ���������������������������������������������������������������������������������������������̋�U����E%�����E�M#M��������   �} tj j �Q�����U�3�t	�E�   ��E�    �M��M��}� uh�aj j1hhaj�%������u̃}� u-��H���    j j1hhahDah�a��?�����   �/�} t�EP�MQ�P�����U���EP�MQ�zP����3���]����������������������������������������������������������������̋�U����EP�M��4���M��$����t2�M��{$������   ~�M��h$��Ph  �UR�PA�����E��h  �EP�M��@$��P� �����E�M�M�M��H���E��]��������������������������������������������̋�U��=�? uh  �EP��!������j �MQ�i9����]�������������̋�U����EP�M��3���M��#����t/�M��#������   ~�M��x#��Pj�UR�c@�����E��j�EP�M��V#��P������E�M�M�M��G���E��]����������������������������������̋�U��=�? uj�EP�� ������j �MQ�%����]����������������̋�U����EP�M��72���M��"����t/�M��"������   ~�M��"��Pj�UR�?�����E��j�EP�M��v"��P�=�����E�M�M�M���F���E��]����������������������������������̋�U��=�? uj�EP� ������j �MQ�q;����]����������������̋�U����EP�M��W1���M���!����t/�M���!������   ~�M��!��Pj�UR�>�����E��j�EP�M��!��P�]�����E�M�M�M���E���E��]����������������������������������̋�U��=�? uj�EP�-������j �MQ�6����]����������������̋�U����EP�M��w0���M��� ����t2�M��� ������   ~�M��� ��Ph�   �UR��=�����E��h�   �EP�M�� ��P�w�����E�M�M�M��E���E��]��������������������������������������������̋�U��=�? uh�   �EP�:������j �MQ�k+����]�������������̋�U����EP�M��/���M�� ����t/�M���������   ~�M�����Pj�UR��<�����E��j�EP�M�����P������E�M�M�M��#D���E��]����������������������������������̋�U��=�? uj�EP�]������j �MQ�/H����]����������������̋�U����EP�M��.���M��'����t/�M��������   ~�M����Pj�UR��;�����E��j�EP�M�����P������E�M�M�M��CC���E��]����������������������������������̋�U��=�? uj�EP�}������j �MQ�9����]����������������̋�U����EP�M���-���M��G����t2�M��;������   ~�M��(��Ph  �UR�;�����E��h  �EP�M�� ��P�������E�M�M�M��]B���E��]��������������������������������������������̋�U��=�? uh  �EP�������j �MQ�w:����]�������������̋�U����EP�M���,���M��W����t2�M��K������   ~�M��8��PhW  �UR� :�����E��hW  �EP�M����P�������E�M�M�M��mA���E��]��������������������������������������������̋�U��=�? uhW  �EP�������j �MQ�7����]�������������̋�U����EP�M���+���M��g����t2�M��[������   ~�M��H��Ph  �UR�09�����E��h  �EP�M�� ��P�������E�M�M�M��}@���E��]��������������������������������������������̋�U��=�? uh  �EP�������j �MQ�/����]�������������̋�U����EP�M���*���M��w����t/�M��k������   ~�M��X��Pj �UR�C8�����E��j �EP�M��6��P�������E�M�M�M��?���E��]����������������������������������̋�U��=�? uj �EP��������j �MQ��6����]����������������̋�U��}�   ���]��������������̋�U��E��]���̋�U��Q�EP�MQ�0������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP�������u�}_t	�E�    ��E�   �E���]�������������̋�U��Q�EP�MQ��6������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP�������u�M��_t	�E�    ��E�   �E���]�������������������������̋�U��E�� ]���̋�U���4�EP�M��(���}   ��   �M������t/�M��������   ~�M�����Pj�UR��5�����E��j�EP�M�����P������Ẽ}� t,�M��������   �E��M��M��=���E��*  ��U�U܍M��=���E��  �M��}��� ���   ~D�M��j��P�M�����   Q�7������t"�U�����   �U��E�E��E� �E�   ��;��� *   �M�M��E� �E�   j�M������BPj�M�Q�U�R�E�Ph   �M�������QR�M�����P�,����$�E�}� u�E�E؍M��0<���E��A�}�u�M��MԍM��<���E��'��U��E���ЉUЍM���;���E���M���;����]����������������������������������������������������������������������������������������������������������������������������̋�U��Q�=�? u$�}A|�}Z�E�� �E���M�M��E���j �UR�������]���������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �O#���E��E��Hp#8t�U��zl ��   j�������E�    �E��Hh�M�U�;8tI�}� t%�E�P�$b��u�}�tj�M�Q�+�����U�8�Bh�8�M�U�R�b�E������   �j�*������	�E��Hh�M�}� u
j �T3�����E�M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E�������!���E��B/���E܋Hh�M��UR��  ���E�E��M;H�  hN  h8bjh   ������E��}� ��  �U܋rh��   �}��E��     �M�Q�UR�������E؃}� ��  �E܋HhQ�$b��u�U܁zhtj�E܋HhQ��)�����U܋E��Bh�M܋QhR�b�E܋Hp���-  �8���  j������E�    �E��H�|?�U��B��?�M��Q��?�E�    �	�E���E�}�}�M�U�E�f�TPf�Mp?���E�    �	�E���E�}�  }�M�M�U�A��0���E�    �	�M���M�}�   }�U�U�E䊊  ��8�׋8R�$b��u�=8tj�8P�(�����M��8�U�R�b�E������   �j��'������(�}��u"�}�tj�E�P�s(�����l6���    ��E�    �E؋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hH�d�    P��$�h3�P�E�d�    �E�    �E�P�M��A!���E�    �l?    �}�u)�l?   ��b�E��E������M��6���E��}�c�}�u)�l?   ��b�E��E������M���5���E��N�4�}�u.�l?   �M��B����Q�U��E������M��5���E���E�E��E������M��5���EЋM�d�    Y��]����������������������������������������������������������������������������̋�U���,�h3ŉE�V�EP�������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0��@;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E����P�M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E���<�UU��B��MM��A����v����U�E�B�M�A   �U�BP��  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��pDf�DJ�ӋMQ�C  ��3��  �����} t!�}��  t�}��  t�UR��b��u����k  �E�P�MQ��b���9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�\  ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=l? t�EP�  ��3�����^�M�3��5����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���  �M��}�w-�U����y
�$��y
�  ��  ��  �	�  �3���]ÍI �y
�y
�y
�y
�y
 ������������������������������������̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U���,�A���E�    �	�M����M��}�   }�UU��E���-��  �׋�]���������������������������������������������������������̋�U���(  �h3ŉE�������P�M�QR��b���-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj ������ j �M�QRh   ������Ph   ������Qh   �U�BPj ������$j �M�QRh   ������Ph   ������Qh   �U�BPj �����$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3��Q/����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��0���M�����H�y t �M�����P�B�E�M��+���E����E�    �M���*���E���M���*����]������������������������������������̋�U��=U uj��0,�����U   3�]����������̋�U��Q�EP�b�M���    t�U���   P�b�M���    t�U���   P�b�M���    t�U���   P�b�M���    t�U���   P�b�E�    �	�M����M��}�m�U����E�|H<t$�M����U�|
P t�E����M�TPR�b�E����M�|L t$�U����E�|T t�M����U�D
TP�b넋M���   �´   R�b��]���������������������������������������������������������������������������������̋�U��Q�} �  �EP�$b�M���    t�U���   P�$b�M���    t�U���   P�$b�M���    t�U���   P�$b�M���    t�U���   P�$b�E�    �	�M����M��}�m�U����E�|H<t$�M����U�|
P t�E����M�TPR�$b�E����M�|L t$�U����E�|T t�M����U�D
TP�$b넋M���   �´   R�$b�E��]������������������������������������������������������������������������������������̋�U��Q�E���    ��   �M���   @!��   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�B�����M���   R�������E���    t4�M���   �: u&j�E���   Q������U���   P�b����j�M���   R������j�E���   Q�������U���    to�E���   �9 uaj�U���   -�   P�����j�M���   ��   R�{����j�E���   ��   Q�a����j�U���   P�M�����M���   @t8�U���   ���    u&�M���   R�#����j�E���   Q������E�    �	�U����U��}���   �E����M�|H<t:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP������M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h�bj h�   hxbj�������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ�����������j�UR��������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�H�����}� t�E�P�N�����}� t�M��9 u�}��t�U�R�*(�����E��]������������������������������������������̋�U��j�h@�h5�d�    P���SVW�h1E�3�P�E�d�    ����E��E��Hp#8t	�U��zl uDj�% �����E�    ��P�M���lQ�6�����E��E������   �j�!�������<���Pl�U�}� u
j �������E�M�d�    Y_^[��]�����������������������������������������������������������̋�U���@�h3ŉE��E�    �E�    �EP�M��/���M�����Pj j j j �MQ�U�R�E�P������ �E��MQ�U�R�"�����E��E���u8�}�u�E�   �M���!���E��j��}�u�E�   �M��!���E��N�:�M���t�E�   �M��!���E��0��U���t�E�   �M��~!���E���E�    �M��j!���E��M�3��$����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�� ����]�������̋�U���@�h3ŉE��E�    �E�    �EP�M�����M��?���Pj j j j�MQ�U�R�E�P�~���� �E��MQ�U�R�������E��E���u8�}�u�E�   �M��f ���E��j��}�u�E�   �M��J ���E��N�:�M���t�E�   �M��, ���E��0��U���t�E�   �M�� ���E���E�    �M������E��M�3��#����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�{����]�������̋�U���@�h3ŉE��E�    �E�    �EP�M��O
���M������Pj j j j �MQ�U�R�E�P����� �E��MQ�U�R�������E��E���u8�}�u�E�   �M������E��j��}�u�E�   �M������E��N�:�M���t�E�   �M�����E��0��U���t�E�   �M�����E���E�    �M�����E��M�3��!����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�+	����]�������̋�U����E�E��M�Q�U�3��} ���E�}� uhj j7h�ij��������u̃}� u0�����    j j7h�ih|ih�������   �$  3�;U��؉E�uhTj j8h�ij�\�������u̃}� u0�u���    j j8h�ih|ihT������   ��  �U� 3��} ����#E��;E��ىM�uh�hj j=h�ij���������u̃}� u0����� "   j j=h�ih|ih�h������"   �J  3��} ���E�}� uh�hj j>h�ij�~�������u̃}� u0����    j j>h�ih|ih�h������   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R��������P�E��P�MQ������3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V� ���M��UR������������0^]������������������������̋�U��Q�E�    �	�E����E��}�-s�M��U;�u�E����7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]��������������������������������������������̋�U��Q�3����E��}� u	�   �������M�3���]�������������������̋�U��Q3��} ���E��}� u!h�.j h�   h0jj�\�������u̃}� u%j h�   h0jhjh�.������   ��P���U� �3���]������������������������������������������̋�U��Q�S����E��}� u	�   ���4����M�3���]�������������������̋�U��Q3��} ���E��}� u!h�.j h�   h0jj�|�������u̃}� u%j h�   h0jh�jh�.������   ������U� �3���]������������������������������������������̋�U��Q�s����E��}� u	�p ���E�����]���������̋�U��Q�C����E��}� u	�t ���E�����]���������̋�U���,�h3ŉE��EP�M�Q� �����U�Rj j���ċMԉ�U؉Pf�M�f�H�������U�B�E�M��U��E�Pj j(hPkh4kh�j�M�Q�UR�EP������P�H�����M�U�Q�E�M�3��@����]���������������������������������������������������̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]����������������������������������������������������������������������������������������������U��WV�u�M�}�����;�v;���  ���   r�=�S tWV����;�^_u�������   u������r)��$�Ж
�Ǻ   ��r����$��
�$���
��$�d�
���
 �
D�
#ъ��F�G�F���G������r���$�Ж
�I #ъ��F���G������r���$�Ж
�#ъ���������r���$�Ж
�I ǖ
��
��
��
��
��
��
��
�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�Ж
����
�
��
�
�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l�
�����$��
�I �Ǻ   ��r��+��$�p�
�$�l�
���
��
̗
�F#шG��������r�����$�l�
�I �F#шG�F���G������r�����$�l�
��F#шG�F�G�F���G�������V�������$�l�
�I  �
(�
0�
8�
@�
H�
P�
c�
�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l�
��|�
��
��
��
�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����?�E��M�����Ƀ��M�uh�lj j*hlj��������u̃}� u+����    j j*hlh�kh�l�������E���E��?�E���]��������������������������������̋�U�졐?]�����SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ����������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����������������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U��W�}3�������ك��E���8t3�����_��������������������̋�U��j�����]���������������̋�U��E��?]�����������������̋�U��Qj��������?P��a�E��MQ��a��?j�������E���]�����������������̋�U��} thlmj jWh�lj��������u�j �q����]���������������������������̋�U�졔?P��a]�������������̋�U��Q��?P��a�E��}� t�MQ�U�����u3���   ��]��������������������������̋�U��   ]����̋�U����S    ]���������������̋�U���V3��} ���E�}� uhnj jHh�mj��������u̃}� u-�5���    j jHh�mh�mhn�W����3��   �}�v����    3��~�} u�E   �URj ��1P��b�E��MQ�URj��1P��b�E��}� u:�}� @  w�M;M�w�x   ��t�U�U��� bP���������
���0�E�^��]����������������������������������������������������������������������������̋�U����E�����j j�E�Pj ��1Q��b��t�}�u	�E�   ��E�    �E���]�������������������������̋�U���V�E�E��} u�MQ��������   �} u�UR�������3��   �E�    �}�w)�} u�E   �EP�MQj ��1R��b�E���EP�t������C	���    3��e�}� u	�=X5 u%�}� t�� bP�#��������	���0�E��1�MQ�%�������u� bP��������������03���J���^��]����������������������������������������������������������������������̋�U��Q�E�����j j ��1P�,b��u�E������E���]�����������������̋�U�������]����̋�U���<�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� uh(3j jih�nj��������u̃}� u.�����    j jih�nhhnh(3�����������  3Ƀ} ���M̃}� uh@nj jnh�nj�U�������u̃}� u.�n���    j jnh�nhhnh@n����������   �E�E��M��A����U��BB   �E�M�H�U�E��M�Qj �UR�E�P��������E��} u�E��Q�M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj �W������EċE���]��������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�C������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�X������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�������]��������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�5�������]������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP���������]����������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�l ������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�* ������]��������������������̋�U��Q�E�E��M�Q�UR�F�������]����������������̋�U��Q�E�E��M�Q�UR�>�������]����������������̋�U��Q�E�E��M�Q�UR�EP���������]������������̋�U��Q�E�E��M�Q�UR�EP��������]������������̋�U��E��=   vhpoj j8h�nj�e�������u̋UR�EPj ������]����������������������������̋�U����EP�M��'����M����   vhpoj jDh�nj���������u̃}�|5�}�   ,�M��l���� ���   �U�Q#E�E�M������E��1�'�M��@�������   �B�#E�E�M�����E���M������]��������������������������������������������������̋�U���(�EP�M��G����}�|6�}�   -�M���������   �E�B#M�M��M�����E��   �M�����P�U�����   R�X�������t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M��5���� �HQ�M��'�����BP�M�Q�U�R�E�Pj�M�����P������ ��u�E�    �M��f���E���M�#M�M؍M��O���E؋�]������������������������������������������������������������������������������̋�U��=�? u�E���A#E��j �UR�EP�I�����]���������������������������U��WV�u�M�}�����;�v;���  ���   r�=�S tWV����;�^_u�_�����   u������r)��$�P�
�Ǻ   ��r����$�d�
�$�`�
��$��
�t�
��
ĩ
#ъ��F�G�F���G������r���$�P�
�I #ъ��F���G������r���$�P�
�#ъ���������r���$�P�
�I G�
4�
,�
$�
�
�
�
�
�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�P�
��`�
h�
t�
��
�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��
�����$���
�I �Ǻ   ��r��+��$��
�$��
� �
$�
L�
�F#шG��������r�����$��
�I �F#шG�F���G������r�����$��
��F#шG�F�G�F���G�������V�������$��
�I ��
��
��
��
��
ȫ
Ы
�
�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��
����
�
�
(�
�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]���������������������������������̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�������������������������������������������̋�U��j�h`�h5�d�    P���SVW�h1E�3�P�E�d�    �e��E�   �E�    �E�P��������u�E�    �E������E��   �M+M�M܋U�R�E�P�4������E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]������������������������������������������������������������������������������̋�U��hy���a��?]���������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e������@x�E�}� t#�E�    �U��E�������   Ëe��E������O����M�d�    Y_^[��]��������������������������������̋�U��Q�����@|�E��}� t�U��������]�������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e衘?P��a�E�}� t#�E�    �U��E�������   Ëe��E������w����M�d�    Y_^[��]��������������������������������������������̋�U��E��?�M��?�U��?�E��?]�����������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    �}t�}u�T  �}t�}t�}t�}t
�}�F  j �������E�    �}t�}u=�=�? u4jh�
��b��u��?   �� b�������0�E�   �E�E̋M̃��M̃}���   �U����
�$�ܴ
��?Q��a�E�}t�UR��a��?�r��?P��a�E�}t�MQ��a��?�L��?R��a�E�}t�EP��a��?�%��?Q��a�E�}t�UR��a��?�E������   �j ������Ã}� t��   ��   �}t�}t�}t��   �����E؃}� u��   �E؁x\p1uLhY  h�pj�2Q�h������EȋU؋EȉB\�}� t�2Qhp1�U؋B\P�#�������j�M؋Q\R�EP�5  ���E��}� u�L�M��Q�U�}t5�E��H;Mu*�U��E�B�M����M��2k��E�P\9U�r��ˋE��   �M�MċUă��Uă}�w�E����
�$��
����x3�t	�E�   ��E�    �E��EЃ}� u!h4pj h�  h�oj���������u̃}� u.�����    j h�  h�oh�oh4p�,�������������M�d�    Y_^[��]Ë�w�
Ĳ
�
��
�
 �I K�
P�
     ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    j �d������E�    �} u�Eܜ?�E܋Q��a�E��E�   ��Eܠ?�U܋P��a�E��E�   �}� t�}�t
�}����M܉�E������   �j � �����Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U���$�
�$��
�EМ?�MЋ�U�E؃��E��  �EР?�MЋ�U�E؃��E���   �EФ?�MЋ�U�E؃��E���   �EШ?�MЋ�U�E؃��E��   ������E��}� u�����  �M��Q\R�EP��  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h4pj h�  h�oj���������u̃}� u1�����    j h�  h�oh�ph4p�0���������4  �E�P��a�E�}�u3��  �}� uj������}� t
j �������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<� 2�M��	�Uԃ��Uԡ 229E�}�M�k��U��B\�D    ���
�����MЉ�E������   ��}� t
j �9�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë���
�
Է
�
��
L�
 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��Q;Ut�E����E��2k�M9M�s�ً2k�U9U�s�E��H;Mu�E���3���]������������������������������������̋�U�졤?P��a]�������������̋�U���\�����d]�����������������̋�U���<�����`]�����������������̋�U��E��?]�����������������̋�U���$V��?P��a�E�3Ƀ} ���M��}� uh�qj jDhpqj�=�������u̃}� u0�V����    j jDhpqh\qh�q�x������   �  �E�     �}� �_  hLG� b�E�}� ut3�t	�E�   ��E�    �U��U�}� uh�pj jPhpqj��������u̃}� u0�����    j jPhpqh\qh�p��������   ��   h�p�M�Q��a�E��}� ��   3�t	�E�   ��E�    �E܉E�}� uh�pj jVhpqj��������u̃}� uD� bP�1������������0j jVhpqh\qh�p�@������ bP��������V�U�R��a�E��T����E��E�Ph�?��b;E�t
�M�Q��bj�UR�U���u�����    ����� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������̋�U��jj �EP�MQ��  ��]���������������������̋�U��jj �EPj ��  ��]�������̋�U��jj �EP�MQ�  ��]���������������������̋�U��jj �EPj �|  ��]�������̋�U��jj �EP�MQ�Z  ��]���������������������̋�U��jj �EPj �,  ��]�������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj ��  ��]��������������������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj �y  ��]��������������������̋�U��jh  �EP�MQ�G  ��]������������������̋�U��jh  �EPj �  ��]��������������������̋�U��jhW  �EP�MQ��  ��]������������������̋�U��jhW  �EPj �  ��]��������������������̋�U��jj�EP�MQ�  ��]���������������������̋�U��jj�EPj �\  ��]�������̋�U��jj �EP�MQ�:  ��]���������������������̋�U��jj �EPj �  ��]�������̋�U��jj �EP�MQ��   ��]���������������������̋�U��jj �EPj �   ��]�������̋�U����EP�M��w����M�������x t8�M�������H�y�  u$jj �UR�EP�i   ���E�M��5����E���E�    �M��!����E��]��������������������������������̋�U��j �EP������]�����������̋�U��j�hx�d�    P���h3�P�E�d�    �EP�M������E�    �M�M�M������P�E�L#Mu;�} t�M����������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M��*����E��M�d�    Y��]��������������������������������������������������������������̋�U����} uh(sj jdh�rj��������u̋M�M��U�R�o������E��E��H��   u$����� 	   �U��B�� �M��A����G  �-�U��B��@t"�v���� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�a����� 9E�t�T�����@9E�u�M�Q��������u�U�R�^������E��H��  ��   �U��E��
+Hy!hrj h�   h�rj�*�������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P��������E��q�}��t!�}��t�M����U������ T�U���E���E��H�� t7jj j �U�R�������E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P�^������E�M�;M�t�U��B�� �M��A�����E%�   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �h3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M������E�    �(����E�3Ƀ} �������������� u!hLvj h  h�uj�Ⱦ������u̃����� uF������    j h  h�uh�uhLv�������ǅ ��������M������� �����  �E�������������Q��@��   ������P�'������������������t-�������t$������������������� T������
ǅ����������H$�����х�uV�������t-�������t$������������������� T������
ǅ����������B$�� ���ȅ�tǅ ���    �
ǅ ���   �� ��������������� u!h�tj h  h�uj�S�������u̃����� uF�i����    j h  h�uh�uh�t������ǅ��������M�����������U  3Ƀ} �������������� u!h(3j h  h�uj�˼������u̃����� uF������    j h  h�uh�uh(3� �����ǅ��������M������������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���g  ������ �Z  �������� |%��������x��������@s���������
ǅ����    ���������������������������`s����������������������������  �������$���
�E�    �M�����P������R����������   ������P�MQ������R�t  ���E��������U���U����������؉�����u!h`tj h�  h�uj��������u̃����� uF�"����    j h�  h�uh�uh`t�A�����ǅ��������M������������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK���������
�$��
�E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP��������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�������Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ��������D�
�$�0�
�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ����������
�$�t�
�U���0  u�E�   �E��M���  tUǅ|���    �UR�i�����f������������Ph   ������Q�U�R��������|�����|��� t�E�   �&�EP�k�����f��x�����x����������E�   �������U��W  �EP�7�������t�����t��� t��t����y u�� �U��E�P�������E��P�M���   t&��t����B�E���t�����+����E��E�   ��E�    ��t����B�E���t�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������l����MQ�d������E��U���  te�}� u�� �E��E�   �M���h�����l�����l�������l�����t��h������t��h�������h����ɋ�h���+M����M��[�}� u	�� �U��E���p�����l�����l�������l�����t��p������t��p�������p����ɋ�p���+E��E��  �MQ��������d������������   3�tǅ����   �
ǅ����    ��������`�����`��� u!htj h�  h�uj��������u̃�`��� uF�,����    j h�  h�uh�uht�K�����ǅ��������M������������  ��  �U��� t��d���f������f����d�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h�sj�Ú�]  R�j������E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���X�����\����M��A���P�E�P�M�Q������R�E�P�M�Q��X���R��P��a�Ѓ��M���   t$�}� u�M������P�U�R��P��a�Ѓ���������gu*�U���   u�M��²��P�E�P��Q��a�Ѓ��U����-u�M���   �M��U����U��E�P��������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�ٻ������H�����L����   �U���   t�EP豻������H�����L����   �M��� tB�U���@t�EP�	���������H�����L�����MQ������������H�����L����=�U���@t�EP����������H�����L�����MQ������3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��M̋Ũ��U̅���@����D���t{�E��RP��D���Q��@���R������0��T����E��RP��D���P��@���Q�������@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �J  ���U�R������P�MQ�U�R�E�P�{  ���M���t$�U���u������P�MQ��<���Rj0��  ���}� ��   �}� ��   ǅ$���    �E���8����M܉�4�����4�����4�������4�������   ��8���f�f������������Pj��(���Q��0���R�(�������$�����8�������8�����$��� u	��0��� uǅ���������*�M�Q������R�EP��0���Q��(���R�z  ���V�����E�P������Q�UR�E�P�M�Q�T  �������� |$�U���t������P�MQ��<���Rj ��  ���}� tj�E�P��������E�    �v���������������M�����������M�3��������]���
��
�
��
��
��
,�
g�
j�
u�
_�
T�
��
��
 �I ��
L�
i�
W�
b�
 ���
��
��
��
N�
�
��
��
 �
��
��
��
��
��
��
   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�8������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A�]��������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��E����U�
�E�f�A�]�������������������̋�U��3�]�������̋�U����E���]��E���]���������̋�S�܃������U�k�l$���   �h3ŉE��C��M��U��U�C��M��U����U��}�w@�E��$���
�E�   �4�E�   �+�E�   �"�E�   ��E�   ��K�   �E�    �}� ��   �U�P�K��Q�U�R�!�������ul�C�E�}�t�}�t�}�t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ�U�R�E�P��p���Q�B�����h��  �U�P� �����ǅl���    �K�9t�=�  u�SR���������l�����l��� u�C�Q�������M�3��������]��[ø�
��
��
��
��
��
��
��
���������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E�}� |,�}�~�}�t���/�M��U��/�y��/�E��o3�t	�E�   ��E�    �U��U��}� uhwj j9h�vj耢������u̃}� u+�����    j j9h�vhtvhw軼���������E���]���������������������������������������������������̋�U��E��/]�����������������̋�U���@�h3ŉE��E�    �u����E��E�    �E�    �E�    �=�? ��   h�w� b�Eԃ}� u3��  h�w�E�P��a�E��}� u3��  �M�Q��a��?h�w�U�R��aP��a��?h�w�E�P��aP��a��?htw�M�Q��a�E��U�R��a��?�=�? thXw�E�P��aP��a��?��?;M�th��?;U�t]��?P��a�EЋ�?Q��a�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W��?;M�t��?R��a�Eȃ}� t�UȉE�}� t*��?;E�t ��?Q��a�Eă}� t
�U�R�UĉE䡸?P��a�E��}� t�MQ�UR�EP�M�Q�U���3��M�3�������]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh0yj jh�xj���������u̃}� u0�����    j jh�xh�xh0y�2������   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E��M���Qh�   �U��R�Y�����3��} ���E��}� uh�Sj jh�xj�.�������u̃}� u0�G����    j jh�xh�xh�S�i������   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E܋M���Qh�   �U��R�`������Px��t3�t	�E�   ��E�    �U؉U�}� uh�wj j h�xj��������u̃}� u0�7����    j j h�xh�xh�w�Y������   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���MԋU���Rh�   �E��P�L������tS��t3�t	�E�   ��E�    �EЉE�}� uh,Sj j*h�xj�
�������u̃}� u-�#���� "   j j*h�xh�xh,S�E������"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�s���U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�b�����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh0yj jh�yj���������u̃}� u0�����    j jh�yh�yh0y�9������   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E�M���Qh�   �U��R�d�����3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���M��U���Rh�   �E��P�������3Ƀ} ���M��}� uh�Sj jh�yj�И������u̃}� u0�����    j jh�yh�yh�S�������   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}�`�����t&�M;MrhtSj j+h�yj�"�������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E܋M���Qh�   �U��R�O������tS��t3�t	�E�   ��E�    �U؉U�}� uh,Sj j>h�yj��������u̃}� u-�&���� "   j j>h�yh�yh,S�H������"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9�s���M���U+U����E+EԋM���Qh�   �U+U��E�LPQ�e�����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���E����E���t��E�+E������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh0yj jh�Sj�ǔ������u̃}� u0�����    j jh�Sh0zh0y�������   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E�M���Qh�   �U��R�)�����3��} ���E��}� uh�Sj jh�Sj���������u̃}� u0�����    j jh�Sh0zh�S�9������   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���M��U���Rh�   �E��P� ������tS��t3�t	�E�   ��E�    �E܉E�}� uh,Sj jh�Sj�ޒ������u̃}� u-������ "   j jh�Sh0zh,S�������"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�s���U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR�6�����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uhpTj jh�yj��������u̃}� u0�'����    j jh�yhHzhpT�I������   �J  �} u\�U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U�E�Ph�   �M��Q�x�����3���  �} ��   �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U��E�Ph�   �M��Q������3҃} �U��}� uh�Sj jh�yj��������u̃}� u0� ����    j jh�yhHzh�S�"������   �#  �M�M��U�U��}�u5�E��M���E���U����U��E���E��t�M����M�t���y�y�����t&�U;UrhtSj j+h�yj�;�������u̋M��U���M���E����E��M���M��t�U����U�t�E���Et�} u�M�� �}� ��   �}�u�UU�B� �P   �?  �E�  �}�tI�}���t@�}v:�M��9�s���U��	�E���E܋M�Qh�   �U��R�s������tS��t3�t	�E�   ��E�    �U؉U�}� uh,Sj j>h�yj�1�������u̃}� u-�J���� "   j j>h�yhHzh,S�l������"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9�s���M���U+U����E+EԋM�Qh�   �U+U��E�LQ苹����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��w����MQ�UR�EP�MQ�M�����P�.   ���E�M��J����E��]�������������������������̋�U����E�    �E��Q�U�j j �EP�MQ��b�E�}� u3���   �}� ~63�u2�����3��u��r#h��  �E�L Q�Ϗ����P�8������E���E�    �U�U��}� u3��s�E�P�M�Q�UR�EP��b��u�H�F�} uj j j j j��M�Qj �U�R��a�E��!j j �EP�MQj��U�Rj �E�P��a�E��M�Q�T������E���]��������������������������������������������������������������������������̋�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�n������.�}���  t%3�u!h�zj h�   h`zj�C�������u̋�]��������������������������̋�U���$�} t�} v	�E�   ��E�    �E�E��}� uh0yj jh`{j�׉������u̃}� u0�����    j jh`{h<{h0y�������   �(  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9�s���U��	�E+E��E�M���Qh�   �U��E�PQ�S�����3���   3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E��M���Qh�   �U��R�������tS��t3�t	�E�   ��E�    �U܉U�}� uh,Sj jlh`{j豆������u̃}� u-�ʩ��� "   j jlh`{h<{h,S�������"   ��   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E�}� v�M����t�E���E�M���M��܋U����:u2�} t!�}s�  j�MQ�UR�EP�V������M���M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E؋M���Qh�   �U��R�������E�    �E�    �E�E��	�M���M�U����t4�M����/t�E����\u�U���U���E����.u�U�U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR�S������E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9�s���M��	�U���UԋE���Ph�   �M��Q�������}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR訢�����}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R�r������   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR�7������}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9�s
���E��	�M(���MЋU���Rh�   �E$��P�������3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9�s���M��	�U���ŰE���Ph�   �M��Q臭�����} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���EȋM���Qh�   �U��R�"������} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9�s
���E��	�M ���MċU���Rh�   �E��P辬�����}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9�s���M��	�U(���U��E���Ph�   �M$��Q�Y�����3҃} �U��}� u!h�|j h�   hH|j�+�������u̃}� u3�D����    j h�   hH|h$|h�|�c������   �   �}� tw3�t	�E�   ��E�    �U��U܃}� u!h�{j h�   hH|j�������u̃}� u0�Ģ���    j h�   hH|h$|h�{�������   �蔢��� "   �"   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���]��������̋�U����} |�}}	�E�   ��E�    �E��E��}� u"h�~j jqh8~j�w}������u��w���}� u.茠���    j jqh8~h~h�~讗��������   �}�t�U���t	�E�    ��E�   �E�E�}� u"h }j jvh8~j��|������u�ww���}� u+�����    j jvh8~h~h }�.���������/�}�u�U��� ��E��� �M��U�E��� �E���]������������������������������������������������������������������������������������������̋�U����} |�}}	�E�   ��E�    �E�E��}� u%h�~j h�   h8~j��{������u�dv���}� u0������    j h�   h8~hh�~������������c�}�u�U�� !�Q�E�� !�M��}�uj��<b�U�� !�'�}�uj��<b�M�� !��U�E�� !�E���]��������������������������������������������������������������̋�U��Q�xS�E��M�xS�E���]������������������̋�U��xS]����̋�U��j�hP�h5�d�    P���PP  ��y���h1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�P�����ƅ���� h�  j ������Q�3�����3�f������h�  j ������P������ƅЯ�� h�  j ��ѯ��Q��������} |�}|����*  �E�    �}��   h� �b����   j h  h8~hx�h�j
h   ��п��R�EP�������P豉����h���b�} t�M�������
ǅ����Ԅ������R��bhȄ��b��п��P��bh(��b�s��ǅ���������=  �} ��   ǅ̯��    �,������ȯ�������     �UR�EPh�  h   ��Я��Q�E�������̯����̯�� }*j h*  h8~hx�hl*j"j�ʛ���R�Wu���� 躛����ȯ�����̯�� }8j h-  h8~hx�h�hJh   ��Я��R������P�s������}uV�} tǅ������
ǅ����܃j h2  h8~hx�h�������Ph   ��п��Q蓜����P������j h4  h8~hx�h����Я��Rh   ��п��P�q����P�݇�����}u�M��� ��t8j h9  h8~hx�hH�h@�h   ��п��P�2q����P萇����j h:  h8~hx�h�h(h   ��п��Q��p����P�X������} ��   ǅį��    �=�����������0����     ��п��P�MQ�URhԁh�  h   ������P�z������į����į�� }*j hA  h8~hx�hl*j"j�ϙ���Q�\s���� 这�����������į�� }8j hD  h8~hx�h@JhJh   ������P�������P�x������:j hH  h8~hx�hh���п��Qh   ������R踚����P�<�����ǅ����    ǅ����    j�������Ph   ������Q������R虌����������j hM  h8~hx�h��j"j������P�kr���� ������ t8j hO  h8~hx�h�h@h   ������Q軙����P蔅�����=�S u�=�S �#  ǅ����    ǅ����    j�ev�����E�   ��S��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un��S��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j蔈����Ã����� �D  �=xS t?ǅ����    ������R������P�MQ�xS����tǅ����   ������������������ ��   �E��� ��t>�U�<� !�t1j ������P������Q�w����P������R�E�� !Q��b�U��� ��t������Q��b�U��� ��twƅп�� �} t9j h�  h8~hx�h�j
h   ��п��Q�UR胏����P�;�������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�������������E������   ��}uh� �$bË������M�d�    Y_^[�M�3��ڙ����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���\�  �o���h1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q������3�f������h�  j ������P�������ƅ���� h�  j ������Q������3�f��Џ��h�  j ��ҏ��P�Û�����} |�}|����.  �E�    �}��   h� �b����   j h�  h8~h��h`�j
h   ��Я��Q�UR�c�����P�}����h ���b�} t�E������
ǅ���؋�����Q��bhċ��b��Я��R��bh����b�i��ǅ���������A  �} ��   ����� ��ȏ��������     �MQ�URh�  h   ��Џ��P�ڈ������̏����̏�� }*j h  h8~h��hl*j"j蠑���Q�-k���� 萑����ȏ�����̏�� }8j h  h8~h��h�h�Nh   ��Џ��P�p�����P�I~�����}uV�} tǅ���Ԋ�
ǅ�����j h  h8~h��h؉�����Qh   ��Я��R������P��}����j h  h8~h��hh���Џ��Ph   ��Я��Q�Zg����P�}�����}u�U��� ��t8j h  h8~h��h�h�h   ��Я��Q�g����P�f}����j h  h8~h��h��h��h   ��Я��R��f����P�.}�����} ��   ǅď��    ����� �����������     ��Я��Q�UR�EPh��h   h   ������Q� �������ď����ď�� }*j h  h8~h��hl*j"j襏���R�2i���� 蕏�����������ď�� }8j h  h8~h��hHOh�Nh   ������R�u�����P�N|�����:j h"  h8~h��h(���Я��Ph   ������Q�9�����P�|����ǅ����    j h(  h8~h��hx�j"jj�������Rh   ������Pj �ב����P�\h���� ������������ t8j h*  h8~h��h��h@�h   ������Q�������P�{�����=�S u�=�S �#  ǅ����    ǅ����    j�Pl�����E�   ��S��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un��S��������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j�~����Ã����� �g  �=xS t?ǅ����    ������R������P�MQ�xS����t������������ǅ����   ������ �  �E��� ���[  �U�<� !��J  �E�� !Q�Db����������t�Jj ������R������P��l����P������Q�U�� !P��b��t��   � b��t��   ǅ���    j h{  h8~h��h��j"jj�������Qh   �����R�����P������P�e���� ���������� t>�����Pt5j ������Q������R�&l������P������P�M�� !R��b�@����� v������������j ������Q�����R�����P�M�� !R��b�E��� ��t������R��b�E��� ��ty3�f��Я���} t9j h�  h8~h��h`�j
h   ��Я��P�MQ��|����P�x������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ�u������������E������   ��}uh� �$bË������M�d�    Y_^[�M�3�袎����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���@�h3ŉE��E�    �m���E��E�    �E�    �E�    �=�? ��   h�w� b�Eԃ}� u3��  h��E�P��a�E��}� u3��  �M�Q��a��?h�w�U�R��aP��a��?h�w�E�P��aP��a��?h��M�Q��a�E��U�R��a��?�=�? thXw�E�P��aP��a��?��?;M�th��?;U�t]��?P��a�EЋ�?Q��a�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W��?;M�t��?R��a�Eȃ}� t�UȉE�}� t*��?;E�t ��?Q��a�Eă}� t
�U�R�UĉE��?P��a�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��-�����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} u3��k  3��} ���E��}� uh��j j7h��j� b������u̃}� u0�9����    j j7h��hh�h���[|�����   �  �} t�U;U��   �EPj �MQ�������3҃} �U��}� uhL�j j=h��j�a������u̃}� u-评���    j j=h��hh�hL���{�����   �~�M;M҃��U�uh�j j>h��j�5a������u̃}� u-�N���� "   j j>h��hh�h��p{�����"   ��   ��MQ�UR�EP�<o����3���]�������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����������������������̋�U���D�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� u!h(3j h�   h0�j��_������u̃}� u1�����    j h�   h0�h�h(3�z��������Z  3Ƀ} ���M̃}� u!h@nj h�   h0�j�l_������u̃}� u1腂���    j h�   h0�h�h@n�y���������   �E�E��M��AB   �U�E�B�M�U��E��@����M�Qj �UR�E�P�3������E��} u�E��   �M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj �hy�����EċE�H���M��U�E��B�}� |!�M�� 3�%�   �E��M����E���M�Qj �y�����E��E���]��������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�u������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ��h������]����������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�m������]������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ��k������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�!h������]��������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP��l������]����������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�k������]��������������������̋�U��Q�E�E��M�Q�UR�d������]����������������̋�U��Q�E�E��M�Q�UR�<^������]����������������̋�U��Q�E�E��M�Q�UR�EP��]������]������������̋�U��Q�E�E��M�Q�UR�EP�u������]������������̋�U��j
j �EP�_����]���������̋�U��EPj
j �MQ�a����]���������������������̋�U��EP�8}����]�������������̋�U��EP�MQ�`c����]���������̋�U��j
j �EP�K�����]���������̋�U��EPj
j �MQ�t����]����������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� ������������������������������������������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ����������������������������XY�$�����������XY�$�����������XY�$����������̋�U���SVWd�5    �u��E�.j �EP�M�Q�UR�*i���E�H����U�Jd�=    �]��;d�    _^[��]� ����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�s���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�gs���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�s���� �E�_^[�E���]��������������������̋�U��E�HQ�U�B(Pj �M�QR�Z����]� �����������������������̋�U����E�    �E�0�h�M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ�Z���E�E�d�    �E��]����������������������������������̋�U��Q��E�H3M�}��j �MQ�U�BP�M�QRj �EP�M�QR�EP��q���� �E��E���]��������������������̋�U���8S�}#  u�.1�M��   ��   �E�    �Eܠ1�h�M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M���a�����   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]��������������������������������������������������������������������̋�U��QS��E�H3M�|���M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ�2p���� �U�z$ u�EP�MQ�_p��j j j j j �U�Rh#  �W�����E��]�c�k ��   [��]���������������������������������������������������̋�U��Q�} �E�HSV�pW�M�����|8����u�uQ���E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v�/Q���M�_��^��[��]��������������������������������̋�U��EV�u���_�����   �N��_�����   ��^]��������������������̋�U���_�����   ��t�M9t�@��u��   ]�3�]�������������������̋�U��V�[_���u;��   u�K_���N���   ^]��:_�����   �x t�H;�t���x u�^]�1P���V�P^]��������������������������U��SVWUj j h(4�u�c��]_^[��]ËL$�A   �   t2�D$�H�3��iy��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h04d�5    �h3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y04u�Q�R9Qu�   �SQ� !�SQ� !�L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������������������̋�U��Q�} t��}��E�P�V  ���M��} t
��  �U���]��������������������������̋�U�����}��E�P�
  ���E��=�S t�]�M�Q��  ��E���E���]�������������������������������̋�U��QV�}���=�S t�E�P�  �����w  ����M�Q�  ��^��]�������������������������������̋�U����} t^��}��E�P��  ���E�M#M�U��#U�ʉM��E�;E�t'�M�Q�Z  ��f�E��m���}��U�R�  ���E��E�M���} t)�=�S t�UR�EP��  ���M��	�U�    �   ��]��������������������������������������������̋�U��E%����P�MQ�
z����]��������������������̋�U�����}��E�P��  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�`  ��f�E��m���}��U�R�  ���E�=�S tB�EP�MQ��  ���E�U�#���E�#��;�t�E�E�   ����E�E����E��]������������������������������������������������̋�U����} 	 u>�}�u8��}��E�%=  ==  u$�=�S t�]��M�����  ���  u�;��7j h[  hX�h4�h���U������R�EPj ��e����P�]������]��������������������������������������̋�U����O��� �E�����F���R	  �}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]�������������������������̋�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]��������������������������������������������������������������������������������������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��������������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�������������������������������������̋�U��Q�yI���E��E�P�)  ����]������������������̋�U��Q�]��e���U��E�P��  ����]��������������̋�U����E%�E�]��M�Q�   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R��  ���E��E�P�;G�����]��M�Q�2   ����]�������������������������������������������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]��������������������������������������������������������������������������������������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]��������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]��������������������������������������������̋�U��Q�E��  �E�P��B������]�������������������̋�U��dS]����̋�U��tS]����̋�U�����O���E��E��Hp����Ƀ��M��U�U��E����E��}�wC�M��$��C�U��Bp���M��Ap�   �U��Bp����M��Ap�   �   �8�����u3�t	�E�   ��E�    �E�E�}� u!hؑj h�   h`�j��B������u̃}� u.��e���    j h�   h`�h0�hؑ�]���������E���]ÐoCjCBCVC�����������������������������������������������������������������������̋�U��j�h��h5�d�    P��SVW�h1E�3�P�E�d�    �=��tAj�C�����E�    h�h��,a�������E������   �j�V����ËM�d�    Y_^[��]�����������������������������������������������̋�U��j�h��h5�d�    P��SVW�h1E�3�P�E�d�    �} ��   j�ZB�����E�    �E�x t.�M�QR�$b��u�E�xtj�M�QR�V�����E������   �j�7U����ËE�8 tcj��A�����E�   �M�R�V^�����E�8 t#�M��: u�E�8�t�M�R�*i�����E������   �j��T����ËE� 𭺋M�A�j�UR�rU�����M�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��EP�A����]�������������̋�U����E�    �} |�}�} u3��  he  hL�jjj�a�����E��}� u�b���    3��  hj  hL�jjh�   �Ta�����M���U��: u j�E�P�ZT�����Sb���    3��8  hp  hL�jjh   �a�����E��M��U��Q�}� u0j�E��Q�T����j�U�R��S������a���    3���   h��E��Q�P  ���UR�EP�M��R�z  ����u3�E��Q�/\�����U��P� g����j�M�Q�S�����E�    �x�U��BP�M���BP�6@������tDj�M��QR�^S�����E��Q��[�����U��P��f����j�M�Q�4S�����E�    ��U��B�    �M��Q�   �E���]���������������������������������������������������������������������������������������������������������������������������������̋�U��VW�} t0�} t*�E;Et"�u�6   �}�M�    �UR�Y����_^]�������������������������������̋�U��EP�MQ�M����]���������̋�U��j�h �h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �(I���E�h�  hL�jjj�^�����E�}� u�_���    3��   ��R���:V���E�M��Ql��E�M��Qh�Pj�q=�����E�    �E�Q�X�����E������   �j�wP�����j�9=�����E�   �U�BP�b�E������   �j�@P����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������̋�U���U��]����̋�U��j�h0�h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �EԉE؃}� u!h��j h&  h`�j��:������u̃}� u0�^���    j h&  h`�h��h���$U����3��  �2G���E��Q���U܋Bp���M܉Ap�E�    h1  hL�jjh�   �}\�����E�}� �  j�;�����E�   �U܋BlP�M�Q��������E�    �   �j�N����Ã}� ��   �UR�EP�M�Q��  ���E��}� ��   �} th<�UR�F>������t
��?   j��:�����E�   �E�P�M܃�lQ�Y�����U�R�SW�����E܋Hp��u$�8��u�E܋HlQh���X�����
  �E�    �   �j��M�������U�R��V�����E�P��a�����E������   ��M܋Qp���E܉PpËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U������   ��!�����   ��!�����   �@%]���������������������̋�U���   �h3ŉE��} tC�} t�EP�MQ�UR�  ����T�����E���M�TH��T�����T����E��|  ǅd���   ǅh���    �} �O  �M���L�'  �E�H��C�  �U�B��_�  �M��`���hԓ��`���R�{1������\�����\��� t"��\���+�`�����X���t��\������;u3���  ǅl���   ���l�������l�����l���N��X���Q��`���R��l���k���@�Q��O������u"��l���k���@�P��:����9�X���u�뚋�\�������\���hГ��\���R�0������X�����X��� u��\������;t3��$  ��l���|j h�  h`�h��h���X���R��\���Ph�   ��p���Q�4����P�HF������X���Ƅp��� ��p���P��l���Q�UR��  ����t��h�������h�����\����X�����`�����`������t��`�������`�����`�������7�����h��� t�MQ��  ����P����
ǅP���    ��P����U��  �EPj j h�   ��p���Q�UR�S�����E��}� ��   ǅl���    ���l�������l�����l���|��l��� tn��l������U�D
HP��p���Q�S9������t;��p���R��l���P�MQ�  ����t��h�������h����
ǅd���    ���h�������h����l�����d��� t�MQ��  ���E��0��h��� t�UR�  ����L����
ǅL���    ��L����E���MQ�  ���E��E��M�3��r[����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �h3ŉE�ǅX���    ǅT���    �?����D�����D����  ��l���ǅH���   �MQ��@���R��L���Ph�   ��p���Q�UR�Q������u3��  �E���M�THR��p���P��6������u�M���U�D
H�a  ��p���P�y6��������T���h�  hL�j��T���Q�-������X�����X��� u3��  �U���E�LH��8����U�E�L���<���j�Uk��E�L$Q��0���R�H@�����E�H��\���j h  h`�h\�hؓ��p���R��T�����P��X�����Q�GV����P��A������X������E���M�TH��L����E�M�T�j��L���R�Ek��M�T$R�?�����}�
  �E��@����H��H�����l����L���T����(�����,���ǅ`���    ���`�������`�����`���;�H�����   �U��`�����l����R;�uJ��`��� t=��`�����l������D���l�����A��`�����l�����(����Ћ�,����L��]�V��`�����l����ЋT���d�����h�����`�����l�����(�������,����T���d�����(�����h�����,����#�����`���;�H�����   j�E�HQ�U�BP��8���Qjh��jj �B���� ����   ǅ$���    ���$�������$�����$���s$��$�����E8������  ��$���f��U8�����h�   �4!P��8���Q��=������u��l����B   ���l����@    ���l����A    ��l����E�H�
�U��l����H���   �}u�U��@����B�MQ�Uk���H��Ѓ���tG�M���U��8����D
Hj��X���Q�"D�����U�E��<����L��U��\����B3��   ��8���<t{�M���U�D
PP�$b��uc3�uj j h[  h`�j�.������u�j�E���M�TPR�C����j�E���M�TTR�C�����E���M�DL    ��X��� t��X����   �E���M��X����TP�E���M�DH�M�3��GU����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�    �E�    �E�    �E�U  ht  hL�j�E�P��'�����E�}� u3��  �M���M��U���U��E��  �M��   �E�   �	�U����U��E����M�THRh�Z�E�k���@�Qj�U�R�E�P�Q&�����}�}kj h�  h`�hȔh��hГ�M�Q�U�R�%����P��;�����E������M�THR�E����M�THR��/������t�E�    �  �}� ��   �E�xP tD�M�QPR�$b��u33�uj j h�  h`�j�O+������u�j�U�BPP�d@�����M�yT tD�U�BTP�$b��u33�uj j h�  h`�j�+������u�j�E�HTQ�@�����U�BT    �E�@L    �M�U�QP�E�M��HH�E���   ��   j�U�R��?�����E�xP tD�M�QPR�$b��u33�uj j h�  h`�j�t*������u�j�U�BPP�?�����M�yT tD�U�BTP�$b��u33�uj j h�  h`�j�'*������u�j�E�HTQ�<?�����U�BT    �E�@L    �M�AP    �U�BH    �E�@h�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����   �h3ŉE��|5���   �E�E��(�E��M�� �M�U��,�U��E�   �E��   �E��E��   �E�    �} u3��-  �} t�} u3��  �M���Cuv�E�H��ukj h�  h`�hL�h��h���UR�EP��L����P�t8�����} t3ɋUf�
3��Mf�A3ҋEf�P�} t	�M�    �E�  �UR�,�����E��}��   s0�EP�M�Q�I,�������  �UR�E�P�1,��������   ǅ@���    ǅD���    �MQ��H���R�U)������t3��  ��H���P�M�Q��H���R��*������u3���   �E��H�U��
��H���P�M�Q�U�R�5-�����E���t�}��   s�U��@����E���D����
ǅ@����j h�  h`�hL�hX���D�����Q��@���R�E�P�M�Q�M%����P�
7�����} tj�U�R�EP�!5�����} tj�M�Q�UR�	5����j h  h`�hL�h���E�P�MQ�UR�#K����P�6�����E��M�3��M����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�]�������̋�U����E�E��E�    �	�M����M��U�;U}A�E����E�j h  h`�h$�hp��M��Q�R�EP�MQ�����P�t5������E�    ��]��������������������������������������������̋�U���h�   j �EP��P�����M���u3���  �E���.uX�U�B��tMj h*  h`�h �h �j�M��Qj�U�   R� #����P�4�����Eƀ�    3��e  �E�    �	�M����M�h��UR�������E��}� u����1  �EE���M��}� uI�}�@sC�U���.t:j h8  h`�h �h(��E�P�MQj@�UR�f"����P�#4�����   �}�uI�}�@sC�E���_t:j h;  h`�h �h8��M�Q�URj@�E��@P�"����P��3�����_�}�uT�}�sN�M���t	�U���,u=j h>  h`�h �h@��E�P�MQj�U�   R�!����P�w3���������)�E���,u��M���u��U��E�L�M����3���]����������������������������������������������������������������������������������������������������������������������������������������̋�U��j hT  h`�hМhH��EP�MQ�UR��F����P�2�����E�H@��t�U��@Rh@�j�EP�MQ������U���   ��t!�M���   Qh��j�UR�EP�P����]����������������������������������������������̋�U����EP�M���0���M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M��'!��P�.   ��$�E�M��E���E��]�������������������������̋�U��� �} ~,�EP�MQ�%  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R��a�E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R�$����P�?�����E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R��a��u
�Y  �T  j j �E�P�M�Q�UR�EP��b�E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR��b��u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�#����P�>�����E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ��b��u�V�T�}  u+j j j j �U�R�E�Pj �M$Q��a�E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P��a�E��}� t�M�Q�@�����U�R�
@�����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U����EP�M��,���M��7����U���   �P�� �  �M�M��A���E��]����������������������������̋�U��j �EP������]�����������̋�U��h  �EP�-����]�������̋�U��h  �EP��,����]�������̋�U��j�EP��,����]����������̋�U��j�EP�,����]����������̋�U��j�EP�,����]����������̋�U��j�EP�g,����]����������̋�U��j�EP�G,����]����������̋�U��j�EP�',����]����������̋�U��h�   �EP�,����]�������̋�U��h�   �EP��+����]�������̋�U��j�EP��+����]����������̋�U��j�EP�+����]����������̋�U��j�EP�+����]����������̋�U��j�EP�g+����]����������̋�U��h  �EP�D+����]�������̋�U��h  �EP�$+����]�������̋�U��hW  �EP�+����]�������̋�U��hW  �EP��*����]�������̋�U��h  �EP��*����]�������̋�U��h  �EP�*����]�������̋�U��j �EP�*����]����������̋�U��j �EP�g*����]����������̋�U���E=�   ���]������������̋�U��Qh  �EP�#*������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP��)������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�)������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�3)������u�M��_t	�E�    ��E�   �E���]��������������������̋�U����EP�M��(���M$Q�U R�EP�MQ�UR�EP�MQ�M��{��P�2   �� �E�M���<���E��]�����������������������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP��a�E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP�J����P�6�����E���E�    �M�M��}� u3��a�U���Rj �E�P��C�����M�Q�U�R�EP�MQj�UR��a�E��}� t�EP�M�Q�U�R�EP��b�E��M�Q��8�����E���]�����������������������������������������������������������������������̋�U��Q�E�x  toj?h��jhd  j�C9�����E��}� u
�   �   �MQ�U�R��   ����t!�E�P�8����j�M�Q�#,�����   �}�U�ǂ�      ��E�@�E���   @tJ�M���   �´   R�$b��u0�E���   ���    hh�j jOh�j�������u̋E�M����   3���]����������������������������������������������������������������̋�U����E�    �E�HB�M��U�BD�E��} u�����  �M�M��E�    �U��Rj1�E�Pj�M�Q�0����E�E�U��Rj2�E�Pj�M�Q�����E�E�U��Rj3�E�Pj�M�Q������E�E�U��Rj4�E�Pj�M�Q������E�E�U��Rj5�E�Pj�M�Q�����E�E�U��Rj6�E�Pj�M�Q�����E�E�URj7�E�Pj�M�Q�m����E�E�U�� Rj*�E�Pj�M�Q�L����E�E�U��$Rj+�E�Pj�M�Q�+����E�E�U��(Rj,�E�Pj�M�Q�
����E�E�U��,Rj-�E�Pj�M�Q������E�E�U��0Rj.�E�Pj�M�Q������E�E�U��4Rj/�E�Pj�M�Q�����E�E�U��Rj0�E�Pj�M�Q�����E�E�U��8RjD�E�Pj�M�Q�e����E�E�U��<RjE�E�Pj�M�Q�D����E�E�U��@RjF�E�Pj�M�Q�#����E�E�U��DRjG�E�Pj�M�Q�����E�E�U��HRjH�E�Pj�M�Q������E�E�U��LRjI�E�Pj�M�Q������E�E�U��PRjJ�E�Pj�M�Q�����E�E�U��TRjK�E�Pj�M�Q�~����E�E�U��XRjL�E�Pj�M�Q�]����E�E�U��\RjM�E�Pj�M�Q�<����E�E�U��`RjN�E�Pj�M�Q�����E�E�U��dRjO�E�Pj�M�Q������E�E�U��hRj8�E�Pj�M�Q������E�E�U��lRj9�E�Pj�M�Q�����E�E�U��pRj:�E�Pj�M�Q�����E�E�U��tRj;�E�Pj�M�Q�v����E�E�U��xRj<�E�Pj�M�Q�U����E�E�U��|Rj=�E�Pj�M�Q�4����E�E�U�   Rj>�E�Pj�M�Q�����E�E�U�   Rj?�E�Pj�M�Q������E�E�U�   Rj@�E�Pj�M�Q������E�E�U�   RjA�E�Pj�M�Q�����E�E�U�   RjB�E�Pj�M�Q�����E�E�U�   RjC�E�Pj�M�Q�\����E�E�U�   Rj(�E�Pj�M�Q�8����E�E�U�   Rj)�E�Pj�M�Q�����E�E�U�    Rj�E�Pj�M�Q������E�E�U�¤   Rj �E�Pj�M�Q������E�E�U�¨   Rh  �E�Pj�M�Q�����E�E�U�°   Rh	  �E�Pj �M�Q�~����E�E�U�E����   �M���   Qj1�U�Rj�E�P�N����E�E�M���   Qj2�U�Rj�E�P�*����E�E�M���   Qj3�U�Rj�E�P�����E�E�M���   Qj4�U�Rj�E�P������E�E�M���   Qj5�U�Rj�E�P�����E�E�M���   Qj6�U�Rj�E�P�����E�E�M���   Qj7�U�Rj�E�P�v����E�E�M���   Qj*�U�Rj�E�P�R����E�E�M���   Qj+�U�Rj�E�P�.����E�E�M���   Qj,�U�Rj�E�P�
����E�E�M���   Qj-�U�Rj�E�P������E�E�M���   Qj.�U�Rj�E�P������E�E�M���   Qj/�U�Rj�E�P�����E�E�M���   Qj0�U�Rj�E�P�z����E�E�M���   QjD�U�Rj�E�P�V����E�E�M���   QjE�U�Rj�E�P�2����E�E�M���   QjF�U�Rj�E�P�����E�E�M���   QjG�U�Rj�E�P������E�E�M��   QjH�U�Rj�E�P������E�E�M��  QjI�U�Rj�E�P�����E�E�M��  QjJ�U�Rj�E�P�~����E�E�M��  QjK�U�Rj�E�P�Z����E�E�M��  QjL�U�Rj�E�P�6����E�E�M��  QjM�U�Rj�E�P�����E�E�M��  QjN�U�Rj�E�P������E�E�M��  QjO�U�Rj�E�P������E�E�M��   Qj8�U�Rj�E�P�����E�E�M��$  Qj9�U�Rj�E�P�����E�E�M��(  Qj:�U�Rj�E�P�^����E�E�M��,  Qj;�U�Rj�E�P�:����E�E�M��0  Qj<�U�Rj�E�P�����E�E�M��4  Qj=�U�Rj�E�P������E�E�M��8  Qj>�U�Rj�E�P������E�E�M��<  Qj?�U�Rj�E�P�����E�E�M��@  Qj@�U�Rj�E�P�����E�E�M��D  QjA�U�Rj�E�P�b����E�E�M��H  QjB�U�Rj�E�P�>����E�E�M��L  QjC�U�Rj�E�P�����E�E�M��P  Qj(�U�Rj�E�P������E�E�M��T  Qj)�U�Rj�E�P������E�E�M��X  Qj�U�Rj�E�P�����E�E�M��\  Qj �U�Rj�E�P�����E�E�M��`  Qh  �U�Rj�E�P�c����E�E�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u�W  j�E�HQ������j�U�BP������j�M�QR������j�E�HQ������j�U�BP�����j�M�QR�����j�E�Q�����j�U�B P�����j�M�Q$R�s����j�E�H(Q�b����j�U�B,P�Q����j�M�Q0R�@����j�E�H4Q�/����j�U�BP�����j�M�Q8R�����j�E�H<Q������j�U�B@P������j�M�QDR������j�E�HHQ������j�U�BLP�����j�M�QPR�����j�E�HTQ�����j�U�BXP�����j�M�Q\R�t����j�E�H`Q�c����j�U�BdP�R����j�M�QhR�A����j�E�HlQ�0����j�U�BpP�����j�M�QtR�����j�E�HxQ������j�U�B|P������j�M���   R������j�E���   Q������j�U���   P�����j�M���   R�����j�E���   Q�����j�U���   P�t����j�M���   R�`����j�E���   Q�L����j�U���   P�8����j�M���   R�$����j�E���   Q�����j�U���   P������j�M���   R������j�E���   Q������j�U���   P������j�M���   R�����j�E���   Q�����j�U���   P�����j�M���   R�p����j�E���   Q�\����j�U���   P�H����j�M���   R�4����j�E���   Q� ����j�U���   P�����j�M���   R������j�E���   Q������j�U���   P������j�M���   R�����j�E���   Q�����j�U��   P�����j�M��  R�����j�E��  Q�l����j�U��  P�X����j�M��  R�D����j�E��  Q�0����j�U��  P�����j�M��  R�����j�E��   Q������j�U��$  P������j�M��(  R������j�E��,  Q�����j�U��0  P�����j�M��4  R�����j�E��8  Q�|����j�U��<  P�h����j�M��@  R�T����j�E��D  Q�@����j�U��H  P�,����j�M��L  R�����j�E��P  Q�����j�U��T  P������j�M��X  R������j�E��\  Q������j�U��`  P�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �E�    �E�E��E�    �M�y u�U�z �  jeh��jjPj� �����E�}� u
�   ��  �E���   �   �}��jqh��jj��������E�}� uj�M�Q�k�����   �z  �U��    �E�x �:  j}h��jj�������E��}� u&j�M�Q�!����j�U�R������   �"  �E��     �M�Q>�U��E�Pj�M�Qj�U�R�����E�E�E��Pj�M�Qj�U�R������E�E�E��Pj�M�Qj�U�R������E�E�E��0Pj�M�Qj�U�R�����E�E�E��4Pj�M�Qj�U�R�����E�E�t0�E�P�����j�M�Q�8����j�U�R�*��������;  �E�HQ�  ���@�E�    �U�@!��M�D!�Q�E�H!�H�U�p!�B0�M�t!�Q4�E��    �}� t	�M��   ��E�    �E�    �E�@!�U���    tA�E���   Q�$b��u-�U���    w!hp�j h�   h��j�/�������u̋M���    t<�U���   P�$b��u(j�M���   R�!����j�E���   Q������U�E����   �M�U쉑�   �E�M䉈�   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�   �E�;@!tj�U�P�>�����M�Q;D!tj�E�HQ������U�B;H!tj�M�QR� �����E�H0;p!tj�U�B0P�������M�Q4;t!tj�E�H4Q������]�����������������������������������������������������̋�U���VW�E�    �E�E��E�    �M�y u�U�z �W  jSh��jjPj�!�����E�}� u
�   ��  jYh��jj�c������E��}� uj�E�P������   ��  �M��    �U�z �d  jeh��jj�������E�}� u&j�E�P�����j�M�Q������   �s  �U��    �E�H8�M��E�    �U��Rj�E�Pj�M�Q������E�E�U��Rj�E�Pj�M�Q�{�����E�E�U��Rj�E�Pj�M�Q�Z�����E�E�U��Rj�E�Pj�M�Q�9�����E�E�U��Rj�E�Pj�M�Q������E�E�U�� RjP�E�Pj�M�Q�������E�E�U��$RjQ�E�Pj�M�Q�������E�E�U��(Rj�E�Pj �M�Q������E�E�U��)Rj�E�Pj �M�Q������E�E�U��*RjT�E�Pj �M�Q�s�����E�E�U��+RjU�E�Pj �M�Q�R�����E�E�U��,RjV�E�Pj �M�Q�1�����E�E�U��-RjW�E�Pj �M�Q������E�E�U��.RjR�E�Pj �M�Q�������E�E�U��/RjS�E�Pj �M�Q�������E�E�U��8Rj�E�Pj�M�Q������E�E�U��<Rj�E�Pj�M�Q������E�E�U��@Rj�E�Pj�M�Q�k�����E�E�U��DRj�E�Pj�M�Q�J�����E�E�U��HRjP�E�Pj�M�Q�)�����E�E�U��LRjQ�E�Pj�M�Q������E�E�t@�U�R�o����j�E�P�
����j�M�Q�
����j�U�R�
�����   �b  �E�HQ�  ����   �@!�}��U���   �M���E���   �U�A�B�M���   �E�J�H�U���   �M�P0�Q0�E���   �U�A4�B4�M��   �}� t	�U��   ��E�    �E�    �E�@!�E���    tA�M���   R�$b��u-�E���    w!hp�j h�   h��j�x�������u̋U���    t<�E���   Q�$b��u(j�U���   P�j	����j�M���   R�V	�����E�M䉈�   �U�E����   �M�U艑�   3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�  �E�H;L!tj�U�BP�������M�Q;P!tj�E�HQ�������U�B;T!tj�M�QR������E�H;X!tj�U�BP������M�Q;\!tj�E�HQ������U�B ;`!tj�M�Q R�a�����E�H$;d!tj�U�B$P�B�����M�Q8;x!tj�E�H8Q�#�����U�B<;|!tj�M�Q<R������E�H@;�!tj�U�B@P�������M�QD;�!tj�E�HDQ�������U�BH;�!tj�M�QHR������E�HL;�!tj�U�BLP�����]�����������������������������������������������������������������������������������������������������������̋�U����i����E��E��Hl�M��U�;�t�E��Hp#8u����E���!��]�����������������������������̋�U�졬!]����̋�U���������E��E��Hl�M��U�;�t�E��Hp#8u����E��U����   ��]�������������������������̋�U��h�!�EP�MQ�h����]��������������������̋�U���<�h3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q�������t	�E�    ��U�R�%�����E�   �Z  �E�P�M�Q��������U�U؋E�HQ�U�R�f������t	�E���E�M�U�A+B9E�}�M�Q�������E�    �E�   ��   �U�E�;Bk�M�Q�U�R�f������E؉E�M�Q+U�UċE�P�M�Q������U�BP�M�Q�������U�B��P�M�Q�u�����E�    �E�   �~�U�E�;|B�M�Q�'�����U܁�   ��U܋E�HQ�U�R�0�����E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�������E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3�������]������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ���������u�U�R�EP�������E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������������������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]��������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P�Z������E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�������E��ȋE���]������������������������������������������������������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]����������������̋�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]����������������������������������̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�����������������������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]������������������������������������������������������������������̋�U��h�!�EP�MQ�����]��������������������̋�U����h3ŉE��E�    �E�H
���  f�M��U�B
% �  f�E�M�Q�U�E�H�M�U����E�j@�M�Q�o�������t�E�   �f�U�f��f�U��E�=�  u�E�   �M�U�Q�E�M��U��E�ЋMf�Q�E��M�3������]��������������������������������������������������������������̋�U���   �h3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h`�j h�   h��j��������u̃}� u0����    j h�   h��h��h`��<�����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$����U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p�����Ī�$����E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h�������$� ��E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�����T��$�H��E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q��������}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�������f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3��;����]Ë�:��������/����g�t��~�l�u���  �֤ͤ�  �˥¥ݥ  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����h3ŉE��P%��`�E��} u�   �} }�M�ىM��&��`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP������눋M�3�������]�����������������������������������������������������������̋�U���L�h3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q������f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R������f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3��w�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]������������������������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]���������������������������̋�U����h3ŉE��EPj j j �MQ�UR�EP�M�Q������� �E�UR�E�P�.������E��}�u	�M���M�E�M�3�������]��������������������������������������̋�U���x�h3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h �h�h��h��j�U��R�������P�]������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h �h�hP�hD�j�U��R�z�����P��������E�@�E�    �   �}�   �uK�}� uEj h�   h �h�h�h�j�M��Q�#�����P�������U�B�E�    �Cj h�   h �h�h��h��j�E��P�������P�b������M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q�������U����?  |f�E�f��f�E��M�Q�U�R�������Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�L�������}� },�E���%�   �E��	�M����M��}� ~�U�R��������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P��������M�Q��������U�R�E�P�������M�Q�������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3��8�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�R�E�Q��������E��}� t0�U��Rj�E�HQ��������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR�l�������]��������������������������������������������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y��������������������������������������������������������������������������������̋�U���8�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh(3j jph�2j�	�������u̃}� u.�"����    j jph�2h��h(3�D���������   3Ƀ} ���MЃ}� uh@nj juh�2j��������u̃}� u.�����    j juh�2h��h@n�����������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P�9������E��} u�E��Q�M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �������EȋE���]������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR������]�������������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h(3j h�  h�2j���������u̃}� u.������    j h�  h�2h̬h(3����������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh��������]������������������̋�U��EP�MQ�URh���W�����]����������������̋�U��EPj �MQhΝ�)�����]������������������̋�U��EP�MQ�URhΝ�������]����������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh(3j jph�2j�	�������u̃}� u.�"����    j jph�2h��h(3�D���������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh@2j jsh�2j��������u̃}� u.�����    j jsh�2h��h@2������������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �~������Eă}��t�E���UU�B� �E��x }�����������]��������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh����������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh���z������E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!hحj h�   h�2j��������u̃}� u1�����    j h�   h�2h��hح�;����������  �} t�} v	�E�   ��E�    �U�U�}� u!h`�j h�   h�2j胿������u̃}� u1�����    j h�   h�2h��h`�����������d  �MQ�UR�EP�MQ�URh���)������E��}� }U�E�  �}�tI�}���t@�}v:�M��9�s���U��	�E���E�M�Qh�   �U��R��������}��uu3�t	�E�   ��E�    �M�M��}� u!h$�j h�   h�2j膾������u̃}� u.����� "   j h�   h�2h��h$�����������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9�s
���E���M����U+щU��E�Ph�   �M��U�D
P��������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�������]���������������̋�U���,�E������E�    3��} ���E�}� u!hحj h  h�2j�̼������u̃}� u1������    j h  h�2h��hح����������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!h`�j h  h�2j�3�������u̃}� u1�L����    j h  h�2h��h`��k���������|  �M;M��   ������U��EP�MQ�UR�E��P�MQh����������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9�s���U���E���M+ȉM�U�Rh�   �E�M�TR�R������v����8"u
�l����M������  �`�X�����U��EP�MQ�UR�EP�MQh���������E��UU�B� �}��u"�}�u�����8"u
�
����M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U��E�Ph�   �M��Q�u������}��uu3�t	�E�   ��E�    �E܉E�}� u!h$�j hB  h�2j�3�������u̃}� u.�L���� "   j hB  h�2h��h$��k�������������z�}�t\�}���tS�U���;UsH�E����M+�9�s���U���E����M+ȉM؋U�Rh�   �E��M�TR�������}� }	�E�������E��EԋEԋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�|�����]�����������̋�U����EPj �MQ�UR�EPhΝ�<������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhΝ��������E��}� }	�E�������U��U��E���]������������������������̋�U��j�hp�h5�d�    P���SVW�h1E�3�P�E�d�    �E������E������}�u!�����     �s���� 	   ��������  �} |�E;�Ss	�E�   ��E�    �MԉM܃}� uh��j jMh �j��������u̃}� u<�I����     ����� 	   j jMh �h�h���#������������C  �E���M������ T�D
������؉E�uhԮj jNh �j�j�������u̃}� u<������     �x���� 	   j jNh �h�hԮ�������������   �UR�s������E�    �E���M������ T�D
��t �MQ�UR�EP�MQ膶�����E��U��F������ 	   �&����     �E������E�����3�uh �j jYh �j菵������u��E������   ��MQ�Ѳ����ËE��U�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��UR��������E�}��u;����� 	   3�u!h �j h�   h �j�l�������u̃������   �UR�E�P�M�Q�U�R��b�E��}��u#� b�E��}� t�E�P�������������>�M���U������ T�L����U���E������ T�L�E��U���]������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �}�u蹼���     �q���� 	   ����  �} |�E;�Ss	�E�   ��E�    �M؉M��}� uh��j jCh�j���������u̃}� u9�J����     ����� 	   j jCh�h�h���$���������/  �E���M������ T�D
������؉E�uhԮj jDh�j�n�������u̃}� u9�Ļ���     �|���� 	   j jDh�h�hԮ����������   �UR�z������E�    �E���M������ T�D
��t�MQ�UR�EP�������E��?����� 	   �4����     �E�����3�uh �j jOh�j褱������u��E������   ��EP������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U�츐<  �����h3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uh�j jmh�j�t�������u̃}� u9�ʹ���     �����    j jmh�h��h�����������
  �E���M������ T�D
$�����E��M���t	�U���uo�E��������E�uh̰j juh�j�ү������u̃}� u9�(����     ������    j juh�h��h̰�����������	  �U���E������ T�T�� tjj j �EP�
������MQ���������td�U���E������ T�T��   tA誻���EԋEԋHl3҃y �U�E�P�M���U������ T�Q��b�E�}� ��  �}� t�U�����  ��b�E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M������ T�|
8 ��   �E���M������ T�D
4P�
�������u!h��j h�   h�j��������u̋U���E������ T�T4�U��EЊ�M��U���E������ T�D8    j�U�R�E�P����������u�  �   �M��R�r���������   �E�+E�M+ȃ�v'j�U�R�E�P�x��������u�O  �MЃ��M��K�U���E������ T�UЊ�T4�E���M������ T�D
8   �E����E���  �j�M�Q�U�R���������u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R��a�Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M������ T�
P��b��t�M�+MM�M��U�;U�}�  �� b�E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M������ T�
P��b��t!�M�;M�}�   �U���U�E����E��� b�E��   �   �M���t	�U���u{�E�P�^��������U�;�u�E����E��� b�E��R�}� tG�E�   �   f�M��U�R���������M�;�u�U����U��E���E��� b�E���t�����  �M���U������ T�L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E������ T�R��b��t �E�E��E�������������+�9M�}��� b�E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U������ T�Q��b��t �U�U��U�������������+�9E�}��� b�E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  ��a��t�����t��� u� b�E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E������ T�R��b��t��p���E���p����� b�E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U������ T�Q��b��t�E�    �U��U��	� b�E�}� ��   �}� t0�}�u�P���� 	   肯���M���U�R�Ȥ��������V�L�E���M������ T�D
��@t�M���u3��%�������    �'����     ������E�+E�M�3��������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} uh(sj j.hx�j詢������u̋�?����?�U�U�j:h<�jh   �������E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������������������������������������������������������̋�U����}�u������ 	   3��   �} |�E;�Ss	�E�   ��E�    �M��M��}� uh��j j(h�j�j�������u̃}� u*����� 	   j j(h�h�h��襻����3���E���M������ T�D
��@��]���������������������������������������������������̋�U���!]����̋�U��Q�=`S u�`S   ��=`S}
�`S   h�   h|�jj�`SP�������@�=@ u?�`S   h�   h|�jj�`SQ�[������@�=@ u
�   �   �E�    �	�U����U��}�}�E����!�M��@�����E�    �	�E����E��}�}f�M����U������� T�<�t8�M����U������� T�<�t�M����U������� T�< u�M���ǁ "�����3���]������������������������������������������������������������������������������������̋�U��舢���00��t趥��j�@Q�0�����]�������������������̋�U��}�!r4�}P$w+�E-�!����P�������M�Q�� �  �E�P��M�� Q��b]�������������������������������̋�U��}}#�E��P薟�����M�Q�� �  �E�P��M�� Q��b]�������������������̋�U��}�!r4�}P$w+�E�H������U�J�E-�!����P�S�������M�� Q��b]�������������������������������̋�U��}}#�E�H������U�J�E��P���������M�� Q��b]�������������������̋�U��Q3��} ���E��}� uhLvj j)hȲj�?�������u̃}� u+�X����    j j)hȲh��hLv�z����������U�B��]�������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E؃}� uh(3j j6hP�j胜������u̃}� u.蜿���    j j6hP�h<�h(3辶��������   �U�U��
����� Pj�(������E�    ������ P�.������E܋E�Pj �MQ�Ү���� P�������E�辮���� P�U�R萻�����E������   �蛮���� Pj�������ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP��������]������������̋�U��Q�E�E��M�Q�UR�EP�ʢ������]������������̋�U��Q�E�E��M�Qj �UR蜢������]��������������̋�U��Q�E�E��M�Q�UR�EP�y�������]������������̋�U��Q�E�E��M�Qj �UR�K�������]��������������̋�U����h��3�9�?���M��} t�h���U���E�    �E���?�E���]������������������������̋�U��h��3�9�?����]��������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uhT�j jJh�j�l�������u̃}� u0腼���    j jJh�hĳhT�觳�����   �\  �UR�M��0����M�谘��� �x ��   �M���   ~C�} t�} v�URj �EP������������ *   � �����M؍M��Լ���E���  �} tw3�;U��؉E�uhTj j]h�j蕘������u̃}� u=讻��� "   j j]h�hĳhT�в�����E�"   �M��_����E��x  �U�E��} t	�M�   �E�    �M��1����E��J  �=  �E�    �U�Rj �EP�MQj�URj �M�舗��� �HQ��a�E��}� t
�}� ��   �}� ��   � b��z��   �} t�} v�URj �EP������3�t	�E�   ��E�    �U��U܃}� uh$�j j{h�j�f�������u̃}� u:����� "   j j{h�hĳh$�衱�����E�"   �M��0����E��L�E���� *   �:�����MȍM������E��*�} t�U�E���E�    �M������E���M��ߺ����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP������]��������������̋�U��� �E������EP�M��Ф���M��P���P�MQ�M��B�������   P�MQ�U�R芠�����E�}� u�E��E���E������M��M�M��z����E��]�����������������������������������������̋�U����E�����j �EP�Ŵ��P�MQ�U�R�������E��}� u�E��E���E������E��]���������������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uh8�j jEh��j��������u̃}� u.蘷���    j jEh��h��h8�躮��������  �MQ�M��E����} �  �M�軓����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M�������E��O  �M����M��U���U뱋E��EԍM��ͷ���E��%  �  �MQ�URj��EPj	�M��1�����QR��a�E��}� t�E����EЍM�肷���E���  � b��zt*艶��� *   3ɋUf�
�E������M��M����E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M�蕒��P�M��R�h�������t@�E��H��u,����� *   3ҋEf��E������M��˶���E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M�������QR��a�E��}� u*蕵��� *   3��Mf��E������M��Y����E��   �U��U��M��C����E��   �   �M�跑��� �x u�MQ�������E��M������E��j�`j j j��URj	�M��}���� �HQ��a�E��}� u!������ *   �E������M��ŵ���E�� ��U����U��M�譵���E���M�蠵����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�UR�EP脙����]�����������������̋�U��=�? uh��EP�MQ�UR�T�������j �EP�MQ�UR�:�����]�����������������������������̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!h�j h�   h��j���������u̃}� u3�ڲ���    j h�   h��h��h���������   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���E��M���Qh�   �U��R�$������} t	�E�     �MQ�M������U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h��j h  h��j迎������u̃}� u@�ر���    j h  h��h��h����������E�   �M�膲���E���  �M������P�E�P�MQ�UR�H������E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���M��U���Rh�   �E��P������������MЍM������E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9�s���M��	�U���U��E���Ph�   �M��Q�T������U�9U����E�u!hP�j h  h��j�(�������u̃}� u=�A���� "   j h  h��h��hP��`������E�"   �M������E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM�贰���Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ臯����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uhpTj jh�xj�G�������u̃}� u0�`����    j jh�xh��hpT肥�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U��E�Ph�   �M��Q譶����3҃} �U��}� uh�Sj jh�xj肊������u̃}� u0蛭���    j jh�xh��h�S轤�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9�s
���E��	�M���M܋U�Rh�   �E��P蹵�����Px��t3�t	�E�   ��E�    �E؉E�}� uh�wj j h�xj�w�������u̃}� u0萬���    j j h�xh��h�w貣�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9�s
���E��	�M���MԋU�Rh�   �E��P諴�����tS��t3�t	�E�   ��E�    �EЉE�}� uh,Sj j*h�xj�i�������u̃}� u-肫��� "   j j*h�xh��h,S褢�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9�s���U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR�ó����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uhj jfh��j��������u̃}� u0�6����    j jfh��h��h�X������   ��  3�;U��؉E�uhx�j jgh��j軅������u̃}� u0�Ԩ���    j jgh��h��hx���������   �  �U� �}�tI�}���t@�}v:�E��9�s���M��	�U���UԋE�Ph�   �M��Q�+�����3҃} ��;U��؉E�uh�j jih��j���������u̃}� u0����� "   j jih��h��h��5������"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uhضj jjh��j�~�������u̃}� u0藧���    j jjh��h��hض蹞�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!h��j h�   h��j�t�������u̃}� u0荦��� "   j h�   h��h��h��謝�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ������]�����������������̋�U��j �EP�MQ�UR�EP�T���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!hj h>  h��j��������u̃}� u3�����    j h>  h��h �h�,������   �,  3�;U���؉E�u!hx�j h?  h��j茀������u̃}� u3襣���    j h?  h��h �hx��Ě�����   ��  �U�� �}��tI�}����t@�}�v:�EЃ�9�s���M��	�UЃ��ŰE�Ph�   �Mԃ�Q�������3҃} ��;U���؉E�u!h�j hA  h��j��������u̃}� u3�ޢ��� "   j hA  h��h �h���������"   ��  �}r�}$w	�E�   ��E�    �UȉU܃}� u!hضj hB  h��j�C������u̃}� u3�\����    j hB  h��h �hض�{������   �{  �E�    �MԉM��} t+�U��-�E����E��M����M��U�ڋE�� �؉U�E�M��M�U3�PR�MQ�UR�+����E�E3�QP�UR�EP�����E�U�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} w�} v�U�;U�r��E�;E�rl�M�� �U�;U���؉E�u!h��j hf  h��j�
~������u̃}� u0�#���� "   j hf  h��h �h���B������"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�B���]����������������̋�U���x�h3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uh�j jfhh�j�|������u̃}� u.�����    j jfhh�h8�h��=���������8  �UR�M��Ȋ���} �.  �M��>{��� �x ��   �M�;Msp�U�=�   ~"讞��� *   �E������M��z����E���  �MM��U���M��E���E��u�M��M��M��D����E��  �U����U�눋E��E��M��#����E��  �  �M��z������   ��   �} v�UR�EP�  ���E�M�Qj �UR�EP�MQ�URj �M��Oz��� �HQ��a�E��}� t3�}� u-�UU��B���u	�M����M��U��U��M�膞���E���  蘝��� *   �E������M��d����E���  ��  �E�Pj �MQ�URj��EPj �M���y����QR��a�E��}� t�}� u�E����E��M������E��j  �}� u� b��zt"����� *   �E������M��ڝ���E��7  �M�;M�  �U�Rj �M��Ay��� ���   Q�U�Rj�EPj �M��$y����QR��a�E�}� t�}� t"蚜��� *   �E������M��f����E���  �}� |�}�v"�l���� *   �E������M��8����E��  �E�E�;Ev�M��M��M������E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M�����E��  벋U���U������E��E��M�蜜���E���   ��   �M��x����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"�i���� *   �E������M��5����E��   �Ũ��U�벋ẺE��M������E��t�j�M�Qj j j j��URj �M��|w��� �HQ��a�E��}� t�}� t����� *   �E������M�辛���E���U����U��M�訛���E���M�蛛���M�3��������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�������������������������������������̋�U��EP�MQ�UR�EP�%�����]�����������������̋�U��j �EP�MQ�UR�������]�������������������̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!hX�j h@  hh�j�u������u̃}� u3�����    j h@  hh�h4�hX��9������   �  �} tU�U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U��E�Ph�   �M��Q�h������} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h��j hL  hh�j�t������u̃}� u3�(����    j hL  hh�h4�h���G������   �  �MQ�U�R�EP�MQ�;������E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9�s���M��	�U���U؋E�Ph�   �M��Q�U������y���� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9�s
���E��	�M���MԋU�Rh�   �E��P�̞�����M9M���ډU�u!h �j hd  hh�j�r������u̃}� u0躕��� "   j hd  hh�h4�h ��ٌ�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h(3j h�   h0�j��p������u̃}� u1������    j h�   h0�h �h(3����������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h@2j h�   h0�j�fp������u̃}� u1�����    j h�   h0�h �h@2螊��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �I������Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj ��������E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh���x}�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh���}�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!hحj h  h0�j�Sm������u̃}� u1�l����    j h  h0�h��hح苇���������  �} t�} v	�E�   ��E�    �U�U�}� u!h��j h  h0�j��l������u̃}� u1�����    j h  h0�h��h������������j  �MQ�UR�EP�MQ�URh����{�����E��}� }X3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���M�U���Rh�   �E��P�������}��uu3�t	�E�   ��E�    �U�U��}� u!h$�j h  h0�j��k������u̃}� u.����� "   j h  h0�h��h$�����������m�}� |d�}�t^�}���tU�M���;MsJ�U����E+�9�s���M���U����E+E��M���Qh�   �U��E�LPQ�0������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�
v����]���������������̋�U���,�E������E�    3��} ���E�}� u!hحj h9  h0�j�j������u̃}� u1�5����    j h9  h0�h �hح�T���������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!h��j h?  h0�j�i������u̃}� u1蜌���    j h?  h0�h �h��軃��������  �M;M��   �_�����U��EP�MQ�UR�E��P�MQh���\x�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9�s���U���E���M+ȉM�U���Rh�   �E�M�TAR蜔����������8"u
趋���M�������  �c袋����U��EP�MQ�UR�EP�MQh���w�����E�3ҋE�Mf�TA��}��u"�}�u�[����8"u
�Q����U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�s
���E��	�M���M��U���Rh�   �E��P蹓�����}��ux3�t	�E�   ��E�    �U܉U�}� u!h$�j hf  h0�j�wg������u̃}� u1萊��� "   j hf  h0�h �h$�证��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9�s���M���U����E+E؋M���Qh�   �U��E�LPQ�Ғ�����}� }	�E�������U��UԋEԋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�"v����]�����������̋�U����EPj �MQ�UR�EPh���t�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh���Vt�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uhj jfh��j�-d������u̃}� u0�F����    j jfh��hH�h�h~�����   �  3�;U��؉E�uhx�j jgh��j��c������u̃}� u0�����    j jgh��hH�hx��~�����   �  3ҋEf��}�tK�}���tB�}v<�M��9�s���U��	�E���EԋM���Qh�   �U��R�7�����3��} ����;E��ىM�uh�j jih��j�c������u̃}� u0����� "   j jih��hH�h��A}�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uhضj jjh��j�b������u̃}� u0装���    j jjh��hH�hض��|�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!h��j h�   h��j�wa������u̃}� u0萄��� "   j h�   h��hH�h���{�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�e�����]�����������������̋�U��j �EP�MQ�UR�EP�4���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!hj h>  h��j��^������u̃}� u3������    j h>  h��hX�h�y�����   �A  3�;U���؉E�u!hx�j h?  h��j�|^������u̃}� u3蕁���    j h?  h��hX�hx��x�����   ��  3ҋE�f��}��tK�}����tB�}�v<�MЃ�9�s���U��	�EЃ��E̋M���Qh�   �Uԃ�R������3��} ����;E���ىM�u!h�j hA  h��j�]������u̃}� u3�ʀ��� "   j hA  h��hX�h���w�����"   �  �}r�}$w	�E�   ��E�    �EȉE܃}� u!hضj hB  h��j�/]������u̃}� u3�H����    j hB  h��hX�hض�gw�����   �  �E�    �UԉU��} t0�-   �M�f��U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ�����E�U3�PR�MQ�UR��}���E�U�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} w�} v�M�;M�r��U�;U�rn3��M�f��U�;U���؉E�u!h��j hf  h��j��[������u̃}� u0���� "   j hf  h��hX�h���%v�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�"���]����������������̋�U����  �h3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���h���E�    ��|���E�3Ƀ} �������������� u!hLvj h  h�uj�Y������u̃����� uF�|���    j h  h�uhp�hLv��s����ǅ<��������M��Y}����<����  3��} �������������� u!h(3j h  h�uj�Y������u̃����� uF�&|���    j h  h�uhp�h(3�Es����ǅ8��������M���|����8����!  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U����  ������ ��  �������� |%��������x��������@s����,����
ǅ,���    ��,������������������������`s����������������(�����(����*  ��(����$��;�E�   ������Q�UR������P�h  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ��������$�����$����� ��$�����$���wL��$�����,<�$�<�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR� w�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�v�����Ẽ}� }�E�������M�k�
�������DЉE��  �������� ����� �����I�� ����� ���.�  �� �����T<�$�@<�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  ��������<�$��<�M���0  u	�U��� �U��E�   �EP��t����f�������M��� tW���������   ������ƅ���� �M��.T��P�M��%T��� ���   Q������R������P�Vu������}�E�   �f������f�������������U��E�   �  �EP�Ht���������������� t�������y u�� �U��E�P�X�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ����������������MQ�xs�����E��U��� ��   �}� u�� �E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M��R��P�������Q�rT������t������������������������������d�}� u	�� �M��E�   �U���|�������������������������t��|������t��|�������|����ɋ�|���+U����U��  �EP�rr������x�����d������   3�tǅ���   �
ǅ���    �������t�����t��� u!htj h�  h�uj�R������u̃�t��� uF�u���    j h�  h�uhp�ht�8l����ǅ4��������M���u����4����  ��  �M��� t��x���f������f����x�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h�sj�Ḿ�]  Q�VL�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��.P��P�U�R�E�P������Q�U�R�E�P��h���Q��R��a�Ѓ��E�%�   t%�}� u�M���O��P�M�Q��R��a�Ѓ���������gu)�M���   u�M��O��P�U�R��P��a�Ѓ��M����-u�E�   �E��M����M��U�R��S�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ��X������X�����\����   �U���   t�EP�X������X�����\����   �M��� tB�U���@t�EP��n��������X�����\�����MQ��n���������X�����\����=�U���@t�EP�n�������X�����\�����MQ�n����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R��p����0��d����E��RP��T���P��P���Q��n����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �]  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��+K��P�M��"K������   R��H���P������Q�Sl������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��L���Rj �  ���}� tj�E�P��_�����E�    �"�����������0����M��n����0����M�3���q����]Ð�.�./y/�/�/0P1R/]/G/</k/t/ �I �041R0?1K1 �
5�1�2�6=2"5�1�647�6�2�6�6�9   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�`�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U���@�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h(3j h�   h0�j�FC������u̃}� u1�_f���    j h�   h0�h��h(3�~]��������V  3Ƀ} ���MЃ}� u!h@nj h�   h0�j��B������u̃}� u1��e���    j h�   h0�h��h@n�]���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P�f�����E��} u�E��   �M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj ��\�����EȋE��H���MċU��EĉB�}� |!�M��� 3�%�   �E��M�����E����M�Qj �\�����E��E���]��������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�_����]�������������������̋�U��EP�MQ�UR�EP�s_����]�����������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h(3j h�  h0�j�v@������u̃}� u.�c���    j h�  h0�h��h(3�Z��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh���X����]������������������̋�U��EP�MQ�URh���gX����]����������������̋�U��EPj �MQh���9X����]������������������̋�U��EP�MQ�URh���X����]����������������̋�U��=�? uj �EP�MQ�URh��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h��d�    P��H�h3�P�E�d�    �EP�M��xM���E�    �} t�M�U�3��} ���Ẽ}� uh̼j j^hX�j�->������u̃}� uD�Fa���    j j^hX�hD�h̼�hX�����E�    �E������M���a���E��  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uh�j j_hX�j�=������u̃}� uD�`���    j j_hX�hD�h���W�����E�    �E������M��Za���E��v  �M�M��E�    �U���E�M����M��M��<����t0�M��<������   ~�M��<��Pj�E�P�Y�����E��j�M�Q�M��r<��P�98�����E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} |�}t�}$~.�} t�U�E��E�    �E������M��O`���E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M����M��U���E�M����M�����3��u�E�j�U�R�M���:��P�6������t�E��0�E��Qh  �M�Q�M���:��P�6������t0�U��a|�E��z�M�� �M���U�U��E���7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M���U�E����E��!����M����M��U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4�`]��� "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U���E��t�M��ىMЋUЉU��E������M���]���E��M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U��=�? uj�EP�MQ�URh���������j�EP�MQ�URj �n�����]�������������������������̋�U��j�EP�MQ�UR�EP�4�����]���������������̋�U��=�? uj �EP�MQ�URh��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�hػd�    P��lVW�h3�P�E�d�    �EP�M��6F���E�    �} t�M�U�3��} ���E��}� uh̼j j^h �j��6������u̃}� uN�Z���    j j^h �h�h̼�&Q�����E�    �E�    �E������M��Z���E��U��<  �} t�}|�}$~	�E�    ��E�   �U��U��}� uh�j j_h �j�K6������u̃}� uN�dY���    j j_h �h�h��P�����E�    �E�    �E������M��Z���E��U��  �M�M��E�    �E�    �U���E�M����M��M��X5����t0�M��L5������   ~�M��95��Pj�E�P�#R�����E��j�M�Q�M��5��P��0�����E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E����E��M���U�E����E��E�RPj�j��V���E�U�j�M�Q�M��4��P��/������t�U��0�U��Th  �E�P�M���3��P�/������t0�M��a|�U��z�E�� �E���M�M��U���7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u^�U�;U�uV�u�3��E�RPj�j��BW���u��}��E��U��E�;E�w.r�M�;M�w$�E�RP�U�R�E�P�3���M�3��։EĉU���U���U�} u��E���M�U����U�������E����E��M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�V��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M���U��t�E��؋Mȃ� �ىEĉMȋUĉU��EȉE��E������M��fV���E��U��M�d�    Y_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�t�����]���������������̋�U��=�? uj�EP�MQ�URh��:�������j�EP�MQ�URj ������]�������������������������̋�U��j�EP�MQ�UR�EP�������]���������������̋�U����<����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR�J3�����   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�i   �� �   ��]���������������������������������������������������������������������������������������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}���+���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  �Y:�����    u��  �F:�����   �E�8:�����   �M�E�j�UR�h.������t��++���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u��*����9�����    ty�9�����   �E��9��ǀ�       �M�Q�UR��  ������t�C�M�Q�  ���Ѕ�t+j�EP�+K����hx��M��B=��h0��M�Q�:����/���U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP��C�����E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q�)C������u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�  ��,�	���D���������M��tj�UR�wI�����E�����   �M��������!���   �E�x ��   �M�QR�EP��  ���ȅ���   �`7�����   �U��R7�����   �E��D7���M���   �67���U���   �}$ u�EP�MQ�F����UR�E$P�~F��j��MQ�UR�EP�.�����M�QR�C  ����6���M���   ��6���U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP�  �� ���,���6�����    u��'����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M��EP�M���C���M�����E���]� ��������̋�U��Q�M��E�� ���M��L����]������������������̋�U��Q�M��M��p?���E��t�M�Q�*�����E���]� �����������������̋�U��Q�M��EP�M���G���M�����E���]� ��������̋�U���V�E�8  �u�c  �X4�����    tW�J4�����`0��9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�*������t��   �M�y t��%���U�R�E�P�MQ�U R�EP��>�����E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������������������������������������������������������������������������������������������������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�*������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����������������������������������������������������̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@�l1��ǀ�       ��'���X1�����    ~�J1���   �E�M����E�3��3���]�������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E��0���   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}��v!���M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R�f'���E�    ��E�P�>����Ëe��E�    �M��M��f����E������   �)��/�����    ~��/���   �EԋUԋ���MԉËU�;Uu�� ���E�M�H�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����E�E��}  t�M Q�UR�E�P�MQ�;F�����}, u�UR�EP�Z>����MQ�U,R�K>���E$�Q�UR�EP�M�Q��%�����U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�T   ���E��}� t�EP�M�Q�N����]�������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R�+�����E���-�����   �E���-�����   �M��-���U���   �-���M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP�>�����E��E�    ��   �M�Q�N  ��Ëe��H-��ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�#�����E�    �E�    �E������E�    �   �   �M�U��Q��E�P� 2�����D,���Mȉ��   �6,���Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP�\/������t�M�Q�UR�=����ËEЋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u�*��ǀ     �   ��3���]�����������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR�������t9j�E�P�w"������t'�M��U�B��M��Q�U��P�uF�����M�������@  �U���txj�M�QR�������tYj�E�P�"������tG�M�QR�E�HQ�U�R�*�����E�xu"�M��9 t�U��R�E��Q��E�����U�������   �E�x uZj�M�QR�(������t>j�E�P�!������t,�M�QR�E��P�M�QR�E����P�E�P�)���������[j�M�QR��������tAj�E�P�:!������t/�M�QR�56������t�E���t	�E�   ��E�   ��R���E�������   Ëe�����E������E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�h5�d�    P���SVW�h1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ��5�����E��}�t�}�t+�R�U��R�E�HQ�C����P�U�BP�M�Q��,���)j�U��R�E�HQ�C����P�U�BP�M�Q�R���E�������   Ëe������E������M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h8�h5�d�    P��SVW�h1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR�dD���E�������E�����Ëe������E������M�d�    Y_^[��]�������������������������������������������������̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]������������������������̋�U����$��3Ƀ��    ����]������̋�U���(�} u3���  �E��M��} t�U�B����   �M��9MOC�t�U��:RCC�t�E��@uz�M��9csm�uK�U��zuB�E��x �t�M��y!�t�U��z"�u�E��x u� $�����    u3��I  �$���   �E܋M܋���E܉�   �%  �M��9csm��  �U��z�  �E��x �t�M��y!�t�U��z"���   �E��x u#�#�����    u3���   �#�����   �M��U�U�E�E��M���   ��M��U��B�H���M�U��B�H��U���E����E��M���M�}� ~d�U��E��M��QR�E�P�M�Q�.������t?�#���   �E؋U؋���M؉�} t�U�R�E�P�MQ�U�R�:�����   ��3���]�����������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E��M����M�U���U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u�!�����   �E��M��QR�E�P�������E��!���M􋐈   ��!���M����   ��w!���M����   ��U�������E�� �����U!���   �E�M����E��;!�����    }�-!��ǀ�       �   ��]������������������������������������������������������������������������������������̋�U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!�f ���   �E��U�����M���   �3���]����������������������������������������������̋�U����E�E��M����M�U���U��E�8��G  �M�Q�%�����} ��   �������   �:csm�u~������   �xum������   �y �t(������   �z!�t������   �x"�u1�o�����   �QR��"������tj�R�����   P�1�����>�����   �9csm�um�+�����   �zu\������   �x �t(������   �y!�t�������   �z"�u �} t�����   �E��E�����U��
����M����   ����M�����   ��]���������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U��j�hX�h5�d�    P��SVW�h1E�3�P�E�d�    �e��E�    �M�U�E�������E�P��+����Ëe��E������M�d�    Y_^[��]��������������������������������������������̋�U��j�hx�h5�d�    P��SVW�h1E�3�P�E�d�    �e��E�    �EP�U���E�������M�Q�4+����Ëe��E������M�d�    Y_^[��]����������������������������������������̋�U��j�h��h5�d�    P��SVW�h1E�3�P�E�d�    �e��E�    �EP�U�E�������M�Q�*����Ëe��E������M�d�    Y_^[��]�������������������������������������������̋�U��j�h��h5�d�    P��SVW�h1E�3�P�E�d�    �e��E�    �EP�MQ�UR�EP�U�E�������M�Q��)����Ëe��E������M�d�    Y_^[��]�����������������������������������������������̋�U����} t�����} u�����E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR�&������t�E���뀊E��]������������������������������������������������������������̋�U��j�h �d�    PQSVW�h3�P�E�d�    �e��v�����    u�����E�    ����$�S���M���   j j �	���E�������x��E���������M�d�    Y_^[��]������������������������������������������������̋�U��Q�E�    �	�E����E��M�U�;}'h�$�E����M�Q�L�K-������t����2���]���������������������������������̋�U����} t��z
���E��M�}� t��e
���U�:csm�u/�E�xu&�M�y �t�U�z!�t�E�x"�u��&
���M�Q�B���E��M�Q�B��M���U����U��E����E��}� ~0�M���U��E��H��Q�M�,&��P�������u�   ��3���]�����������������������������������������������������������U���SQ�E���E��EU�u�M�m�� ��VW��_^��]�MU���   u�   Q����]Y[�� �������������������̋�U���@�h3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �M�y ��  �U�z u+�E��Ph  �M�Q0Rj �E�P�_������t�"  j^hP�jj�\�����E�jbhP�jjh�  ��,�����E�jdhP�jjh�  �,�����E�jfhP�jjh�  �,�����E�jhhP�jjh  �,�����E�}� t�}� t�}� t�}� t�}� u�}  �M��    �U�U��E�    �	�E����E��}�   }�M��U���E����E��ۍM�Q�U�BP��b��u�&  �}�v�  �M܉Mă}�~S�U�U��	�E����E��M����t8�E��H��t-�U���E��	�M����M��U��B9E��M�M�� ���j j �U�BP�Ḿ�   Qh   �U�Rjj ������ ��u�  j �E�HQh�   �Uȁ   Rh�   �E��Ph   �M�QRj � ����$��u�E  j �E�HQh�   �U��   Rh�   �E��Ph   �M�QRj �����$��u�  3��M�f���   �U��B �E��@ �M�Ɓ�    �U�Ƃ�    �}�~]�E�E��	�M����M��U����tB�M��Q��t7�E���M��	�U����U��E��H9M�� �  �E��M�f��A   ���h�   �Ú�   R�E�P�����j�Mȁ�   Q�U�R�s����j�E�   P�M�Q�\�����U���    ��   �E���   Q�$b����   3�uj j h�   hؽj�������u�j�M���   ���   R������j�E���   ��   Q�����j�U���   -�   P�����j�M���   R������E��    �M�UЉ��   �E�   �M���   �Ú��   �E���   �Mȁ��   �U���   �E��   �M���   �U�Eĉ��   j�M�Q�����3���   j�U�R������j�E�P������j�M�Q������j�U�R������j�E�P�������   �   �   �M���    tA�U���   P�$b��u-�M���    w!h��j h�   hؽj�>������u̋Eǀ�       �Mǁ�       ����E���   ����U���   � ��M���   �Uǂ�      3��M�3��-����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��������E��E��Hl�M��U�;�t�E��Hp#8u����E��U����   ��]�������������������������̋�U��Q�} u
�#���E���E����   �U��E���]���������������������̋�U����9���E��E��Hl�M��U�;�t�E��Hp#8u�����E��U��B��]����������������������������̋�U��������E��E��Hl�M��U�;�t�E��Hp#8u����E��U��B��]����������������������������̋�U����y���E��E��Hl�M��U�;�t�E��Hp#8u�'���E��E�����]����������������������������̋�U��3�]��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^���������������������������̋�U��Q�E�    �} u3��S  �}��   �	�E����E��M��9M���   �U���U�E���E�M�Q���t�E�H��U�B�;�t�M�A��U�J�+���   �U�B���t�M�Q��E�H�;�t�U�B��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��X�����	�E����E��M�;Ms>�U���t�M��E�;�t�U��M�+���E���E�M���M�3���]������������������������������������������������������������������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U���(�E�E��M�M��U�U��}��g  �E��$���M�Q�U�R��  ���E�}� t�E�E��s�M���Q�U���R��  ���E�}� t�E�E��F�M���Q�U���R�  ���E�}� t�E�E���M���Q�U���R�  ���E�E�E�M�M�E���   �U�R�E�P�Y  ���E�}� t�M�M��F�U���R�E���P�2  ���E�}� t�M�M���U���R�E���P�  ���E܋M܉M��E��i�U�R�E�P��   ���E�}� t�M�M���U���R�E���P��   ���E؋E��*�M�Q�U�R�   ���3���EP�M�Q�U�R�  ����]Ð�����:��������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��+�P�   ����]�����������������̋�U��} t3��} ���D ��E�E]����������������̋�U����} �R  �EP�MQ�Q	  ���E��}� t�E��O  �U��R�E��P�*	  ���E��}� t�E��(  �M��Q�U��R�	  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�g  ���E��}� t�E��e  �U��R�E��P�@  ���E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$����U��R�E��P��  ���E��}� t�E���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��}  �U��R�E��P�X  ���E��}� t�E��V  �M��Q�U��R�1  ���E��}� t�E��/  �E��P�M��Q�
  ���E��}� t�E��  �U��R�E��P��  ���E��}� t�E���  3���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��  �U��R�E��P�g  ���E��}� t�E��e  �M��Q�U��R�@  ���E��}� t�E��>  �E��P�M��Q�  ���E��}� t�E��  �U��	R�E��	P��  ���E��}� t�E���  �M��Q�U��R��  ���E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�b  ���E��}� t�E��`  �E��P�M��Q�;  ���E��}� t�E��9  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���E��}� t�E���  �E��
P�M��
Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���  �E��P�M��Q�]  ���E��}� t�E��[  �U��R�E��P�6  ���E��}� t�E��4  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���   �U��R�E��P��  ���E��}� t�E��   �M��Q�U��R�  ���E��}� t�E��   �E��P�M��Q�s  ���E��}� t�E��t�U��R�E��P�o������E��}� t�M��M��F�U��R�E��P�H������E��}� t�M��M���U��R�E��P�!������E��M��M�E��3���]Ë���Ɍ�������΍��c�{���ӎ<�T������-�Y�����2�^�Ǌߋ�7������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��;�tK�E�E��M�M�U�R�E�P�������E�}� t�M�M���U���R�E��P�\������E�E��3���]�������������������������������������������̋�U��� �E�E��M�M��U��E��
;��   �U�U��E�E�M�Q�U�R��������E�}� t�E�E��s�M���Q�U��R�������E�}� t�E�E��F�M���Q�U��R�������E�}� t�E�E���M���Q�U��R�n������E��E��E�M�M�E��3���]�����������������������������������������������������������������̋�U����i����   �E��} u�E�P�\  ���  �M��U��E��@�M��A�U��z t#�E��H���t�E���Pjh����  ���M��A    �U��: ��   �E�������   �E��x t�M��Q���t�M�Q�O  ����U�R�	  ���E��x uG�M�Qj@h`��u  ����t0�U��z t�E��H���t�E�P��  ����M�Q�1	  ���0�U��z t�E��H���t�E�P�  ����M�Q�?  ���U��z u3��N  �} t�E�   �E���E�    �M�Q�U�R�U  ���E��}� t!�}���  t�}���  t�E�P��b��u3���   j�M��QR� c��u3���   �} t&�E�M�f�Qf��E�M�f�Qf�P�Ef�M�f�H�} ��   �U�=  u4j h1  h8�h��h��h��j@�MQ�Y����P�� ����� j@�URh  �E��HQ��b��u3��Bj@�U��@Rh  �E��HQ��b��u3��j
j�U�   R�E�P������   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�;Eb�}� t\�E�E�+����E��M��U��P�M�R�2�����E�}� u�E��M�T��E���}� }�M����M�	�U����U��3��}� ����]�����������������������������������̋�U��Q�E�Q�������3҃��E�P�M�QR�������3Ƀ����U�J�E�@    �M�y t	�E�   ��U�P��  ���E��M�U��Qjh���c�E�H��   t�U�B%   t�M�Q��u
�E�@    ��]����������������������������������������������������������̋�U���   �h3ŉE��l����   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q��b��u��|����B    �   �  �E�P��|����QR�I�������r  jx�E�P��|����Q��ҁ������  R��x���P��b��u��|����A    �   �G  �U�R��|����Q��������u:��|����B  ��|����A��|�����x����B��|�����x����Q��   ��|����H����   ��|����z tt��|����HQ�U�R��|����Q�S������uQ��|����B����|����A��|�����x����B��|����R�c�������|���;Au��|�����x����B�E��|����Q��u7��x���P��  ����t$��|����Q����|����P��|�����x����Q��|����H��   ��   ��  jx�U�R��|����H��Ɂ������  Q��x���R��b��u��|����@    �   �  �M�Q��|����P�W�������
  ��|����Q��   ��|����P��|����y t7��|����B   ��|����A��|����z u��|�����x����H�   ��|����z tl��|����Q�
�������|���;BuP��|���Pj��x���Q��  ����t2��|����B   ��|����A��|����z u��|�����x����H�2��|����B   ��|����A��|����z u��|�����x����H�   ��|����z ut��|����x th�M�Q��|����P�������uO��|���Qj ��x���R�C  ����t3��|����H��   ��|����J��|����x u��|�����x����Q��|����@��������M�3������]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�Q������3҃��E�P�M�y t	�E�   ��U�P��  ���E��M�U��Qjhp��c�E�H��u
�U�B    ��]��������������������������������������������̋�U���   �h3ŉE��|����   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q��b��u��|����B    �   �  �E�P��|����R�Z
������u`��|����x u��|���Qj��x���R�y  ����t3��|�����x����H��|�����x����B��|����Q����|����P�   ��|����y ut��|����z th�E�P��|����R��	������uO��|���Pj ��x���Q��  ����t3��|�����x����B��|�����x����Q��|����H����|����J��|����@��������M�3������]� ������������������������������������������������������������������������������������������������������̋�U��E�HQ������3҃��E�PjhР�c�M�Q��u
�E�@    ]��������������������������̋�U���   �h3ŉE������   ��|����EP�B  ����x���jx�M�Q��|����B���%���  P��x���Q��b��u��|����B    �   �s�E�P��|����QR��������uF��x���P��  ����t3��|�����x����Q��|�����x����H��|����B����|����A��|����B��������M�3�������]� ������������������������������������������������������������������̋�U��Q�E�H��  �U�J�c�E��E�M��H�U�E��B��]�������������������������̋�U��Q�} t�E���th���UR�X�������u0j�E�Ph  �M�QR��b��u3��Y�}� u��b�K�Fh���EP��������u"j�M�Qh   �U�BP��b��u3����MQ�������E��E���]��������������������������������������������������������̋�U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E��;�u3���ظ   ��]����������������������̋�U���V�E%�  �ȁ�   �щU�j�E�Ph   �M�Q��b��u3��9�U;U�t,�} t&�E�Q��   �����U�P������;�u3���   ^��]������������������������������������̋�U����E�    �E��M��U��E���E��tM�M���a|�U���f�E���'�E���M���A|�U���F
�E����E��M����U��DЉE�뚋E���]������������������������������������̋�U����E�    �E��M��U���U�E���A|	�M���Z~�U���a|%�E���z�M����M��U��E��M���M���E���]�������������������������̋�U���EP�MQ�������]�������̋�U��Q�E=��  u3��G�M��   }�U��!�P�M#��&�U�Rj�EPj��b��u3�f�M��E��U#�]��������������������������������̋�U���EP�MQ�D�����]�������̋�U����h3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ�j������UR�^������E�P�MQ�;������UR�B������E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR������f�E�f��f�E��؋Mf�U�f�Q
�M�3��K����]����������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����'  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tE�U�;U�u.�E�H��  ����ًU��  �����;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���(  �h3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T����A���ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �������|���3Ƀ} ����0�����0��� u!hLvj h  h�uj��������u̃�0��� uI�����    j h  h�uh��hLv�������ǅ ���������T����Q����� �����7  �E��,�����,����Q��@��   ��,���P���������(�����(����t-��(����t$��(�������(�������� T��\����
ǅ\������\����H$�����х�uV��(����t-��(����t$��(�������(�������� T��X����
ǅX������X����B$�� ���ȅ�tǅT���    �
ǅT���   ��T�����$�����$��� u!h�tj h  h�uj��������u̃�$��� uI�1����    j h  h�uh��h�t�P�����ǅ����������T���������������T6  3Ƀ} ���� ����� ��� u!h(3j h  h�uj��������u̃� ��� uI�����    j h  h�uh��h(3�������ǅ����������T����N�����������5  ǅL���    �E������ǅ@���    ���@�������@�����@����q5  ��@���u������ u�Z5  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Uǅ��������ǅ��������ǅp�������ǅ���������E���G�����G����E���E����1  ��L��� ��1  ��G����� |%��G�����x��G�����������P����
ǅP���    ��P�����H�����H���k�	��8����������8�����8�����  �E���%��  �������u\j
��t���R�EP��������~9��t������$u+��@��� uh@  j ������P�n����ǅ����   �
ǅ����    �������)  j
��t���Q�UR����������������t������E��@��� ��   ������ |#��t������$u������d}ǅL���   �
ǅL���    ��L������������� u!h8�j hQ  h�uj��������u̃���� uI������    j hQ  h�uh��h8��������ǅ����������T����k�����������2  ������;�x���~��������H������x�����H�����H�����x����   ��8�����   3�tǅD���   �
ǅD���    ��D������������� u!h��j h]  h�uj���������u̃���� uI������    j h]  h�uh��h���������ǅ����������T���������������1  ��8�����@�����@�����.  ��@����$� ���@��� u	������t��@���u�������u�.  ǅ����    ��T�������P��G���R�o���������   ��L���P�MQ��G���R�9A  ���E���G����U���U��G�������؉����u!h`tj h�  h�uj��������u̃���� uI�����    j h�  h�uh��h`t�������ǅ����������T����O�����������0  ��L���R�EP��G���Q�@  ���-  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �P-  ��G�����<�����<����� ��<�����<���wi��<�����X��$�@����������������D���������������3���������������"�������   ����������������������,  ��G�����*��  ������ u�EP�"������������^  j
��t���Q�UR�U���������������t������E��@��� ��  ������ |#��t������$u������d}ǅ8���   �
ǅ8���    ��8������������� u!h(�j h�  h�uj�h�������u̃���� uI�~����    j h�  h�uh��h(�������ǅ����������T����&����������.  ������;�x���~��������4������x�����4�����4�����x����������������� uE��������Ǆ����   ����������G������������������������������   ������P��G���Qj��������������P�v���������؉����u!h��j h�  h�uj�1�������u̃���� uI�G����    j h�  h�uh��h���f�����ǅ����������T���������������j-  �\*  �+������������������������Q������������������ }���������������������؉������������k�
��G����DЉ�������)  ǅd���    ��)  ��G�����*��  ������ u�UR�>�������d����^  j
��t���P�MQ�q���������p�����t������U��@��� ��  ��p��� |#��t������$u������d}ǅ0���   �
ǅ0���    ��0������������� u!h��j h�  h�uj��������u̃���� uI�����    j h�  h�uh��h��������ǅ����������T����B����������+  ��p���;�x���~��p�����,������x�����,�����,�����x�����p����������� uE��p�����Ǆ����   ��p�������G�����������p������������������   ������R��G���Pj��p�����������R����������؉� ���u!h �j h�  h�uj�M�������u̃� ��� uI�c����    j h�  h�uh��h �������ǅ����������T��������������*  �x'  �+��p�����������������������P���������d�����d��� }
ǅd����������d���k�
��G����DЉ�d����'  ��G�����(�����(�����I��(�����(���.�B  ��(��������$�l��U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅ8���    �*����"�������� �������������   �������%  ��G�����$�����$�����A��$�����$���7��"  ��$��������$�����������0  u������   ��������������  �_  ǅ����    ������ u�UR�W�����f��<�����  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!h��j h�  h�uj�.�������u̃����� uI�D����    j h�  h�uh��h���c�����ǅ����������T���������������g'  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�c���������؉�����u!h�j h�  h�uj��������u̃����� uI�4����    j h�  h�uh��h��S�����ǅ����������T���������������W&  �   �,��������������������������P�_�����f��<�����<���Qh   ��P���R������P�
����������������� t
ǅl���   �*  ������ u�MQ�O�����f��������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h��j h�  h�uj���������u̃����� uI������    j h�  h�uh��h��������ǅ����������T��������������%  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�����u!hx�j h�  h�uj���������u̃����� uI������    j h�  h�uh��hx��������ǅ����������T��������������$  �j  �,��������������������������R�W�����f��������������P���ǅ����   ��P����������  ������ u�UR��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h��j h�  h�uj��������u̃����� uI�����    j h�  h�uh��h���������ǅ����������T����]�����������"  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�����������؉�����u!h��j h�  h�uj��������u̃����� uI�����    j h�  h�uh��h���������ǅ����������T����M�����������!  �0  �+��������������������������P������������������ t�������y u#�� ������������P��������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������a  ������%0  u��������   ��������d����uǅ���������d������������������������� u�MQ��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h��j h6  h�uj��������u̃����� uI�����    j h6  h�uh��h���������ǅ����������T����]�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�����������؉�����u!h��j h:  h�uj��������u̃����� uI�����    j h:  h�uh��h���������ǅ����������T����M�����������  �0  �+��������������������������R������������������%  tx������ u�� ������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������i������ u�� ����������������������������������������t���������t���������������ɋ�����+������������  ������ u�UR��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h��j h�  h�uj蚿������u̃����� uI�����    j h�  h�uh��h���������ǅ����������T����X�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�����������؉�����u!h��j h�  h�uj芾������u̃����� uI�����    j h�  h�uh��h��������ǅ����������T����H�����������  �+  �+��������������������������P��������������������   3�tǅ���   �
ǅ���    ����������������� u!htj h�  h�uj詽������u̃����� uI�����    j h�  h�uh��ht�������ǅ����������T����g�����������  �J  �������� t������f��L���f����������L����ǅl���   �  ǅh���   ��G����� ��G�����������@��������������  ��@��� ��  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h��j h�  h�uj�w�������u̃����� uI�����    j h�  h�uh��h��������ǅ����������T����5����������  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�����u!h0�j h�  h�uj�t�������u̃����� uI�����    j h�  h�uh��h0�������ǅ����������T����2����������  �  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��G�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Zh�  h�sj��d�����]  R������������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�U���U�E�H��P��������������  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!h��j h  h�uj�˹������u̃����� uI������    j h  h�uh��h��� �����ǅ����������T��������������  ��@���t!h��j h  h�uj�O�������u̋����������������������������������������H��P���������������T���蕸��P��h���P��d���Q��G���R��P���P������Q������R��P��a�Ѓ���������   t-��d��� u$��T����6���P������R��P��a�Ѓ���G�����gu3��������   u%��T��������P������P��Q��a�Ѓ����������-u!��������   ��������������������������P��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ��������   t ƅ����0��4�����Q������ǅ����   �*ǅ����   ��������   t��������   ������������% �  �#  ������ u�MQ��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u!h��j h�  h�uj���������u̃�l��� uI������    j h�  h�uh��h���������ǅ����������T���������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�����������؉�h���u!hH�j h�  h�uj豵������u̃�h��� uI������    j h�  h�uh��hH��������ǅ����������T����o�����������  �R  �1����������������d�����d���R躾������x�����|�����
  ������%   �#  ������ u�MQ胾������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������`�����`��� u!h��j h�  h�uj荴������u̃�`��� uI�����    j h�  h�uh��h���������ǅ����������T����K�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�¿��������؉�\���u!h��j h�  h�uj�}�������u̃�\��� uI�����    j h�  h�uh��h��������ǅ����������T����;����������  �  �1����������������X�����X���R膼������x�����|�����  �������� �a  ��������@�'  ������ u�UR�����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������T�����T��� u!h��j h�  h�uj�J�������u̃�T��� uI�`����    j h�  h�uh��h��������ǅ����������T��������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�P���u!hx�j h�  h�uj�:�������u̃�P��� uI�P����    j h�  h�uh��hx��o�����ǅ����������T���������������s  ��  �3����������������L�����L���P�����������x�����|����&  ������ u!�MQ�����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������H�����H��� u!h��j h�  h�uj�!�������u̃�H��� uI�7����    j h�  h�uh��h���V�����ǅ����������T���������������Z  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�V���������؉�D���u!hx�j h�  h�uj��������u̃�D��� uI�'����    j h�  h�uh��hx��F�����ǅ����������T���������������J  �  �5����������������@�����@���R�����������x�����|����V  ��������@�%  ������ u�MQ�f��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������<�����<��� u!h��j h  h�uj��������u̃�<��� uI� ����    j h  h�uh��h��������ǅ����������T��������������#  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�8���u!hx�j h  h�uj�ڬ������u̃�8��� uI������    j h  h�uh��hx�������ǅ|���������T���������|����
  �{  �2����������������4�����4���R�h��������x�����|����"  ������ u�EP�A�����3ɉ�x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������0�����0��� u!h��j h0  h�uj�ī������u̃�0��� uI������    j h0  h�uh��h���������ǅx���������T���������x�����  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�����������؉�,���u!hx�j h4  h�uj贪������u̃�,��� uI������    j h4  h�uh��hx��������ǅt���������T����r�����t�����  �U  �3����������������(�����(���R�B�����3ɉ�x�����|�����������@tG��|��� >|	��x��� s3��x����؋�|����� �ى�p�����t�����������   ���������x�����p�����|�����t����������� �  u(������%   u��p�����t����� ��p�����t�����d��� }ǅd���   �%�����������������d���   ~
ǅd���   ��p����t���u
ǅ����    ��O�����������d�����d�������d�������p����t�����   �������RP��t���P��p���Q�\�����0�������������RP��t���R��p���P�4�����p�����t���������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�s  ��l��� �B  ��������@t[��������   tƅ����-ǅ����   �:��������tƅ����+ǅ����   ���������tƅ���� ǅ����   ������+�����+�������$�����������u��L���Q�UR��$���Pj �m  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��$���Qj0�  �������� ��   ������ ��   ǅ���    �������� �����������������������������������   �� ���f�f������������Rj�����P�����Q�������������� ������� �������� u	����� uǅL��������-��|���P��L���Q�UR�����P�����Q�  ���S����(��|���R��L���P�MQ������R������P�P  ����L��� |'��������t��L���R�EP��$���Qj ��  �������� tj������R论����ǅ����    ������8��� t��8���tǅ����    �
ǅ����   ���������������� u!h(�j h�  h�uj��������u̃���� uI�1����    j h�  h�uh��h(��P�����ǅp���������T����������p����T  �������%  ��@��� �  ǅ����    ���������������������;�x�����  �����������������������������������������  �������$�$����������E�������MQ�0������  ���������E�������MQ迻�����_  ���������E�������MQ��������;  ���������E�������MQ�?������  ���������E�������MQ��������   ���������E�������MQ�|�������   ���������E�������MQ��������h�����l����   3�tǅ����   �
ǅ����    ���������������� u!h��j h.	  h�uj��������u̃���� uF�����    j h.	  h�uh��h��� �����ǅd���������T���������d����'������s�����L�����`�����T���������`����M�3�������]Ë�8�f���J��.��`��#���6�E� �I i�9�-�J�[� �m������h�����~�m����;�����}�   	
B�f���������J���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP��������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U���<  �h3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��&����E�    �8����E�3Ƀ} �������������� u!hLvj h  h�uj�؏������u̃����� uF�����    j h  h�uht�hLv������ǅ��������M�虳��������#  �E�������������Q��@��   ������P�7������������������t-�������t$������������������� T�������
ǅ������������H$�����х�uV�������t-�������t$������������������� T�������
ǅ������������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h�tj h  h�uj�c�������u̃����� uF�y����    j h  h�uht�h�t蘨����ǅ��������M��$���������  3Ƀ} �������������� u!h(3j h  h�uj�ۍ������u̃����� uF�����    j h  h�uht�h(3������ǅ��������M�蜱��������&  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���  ������ �	  �������� |%��������x�������������������
ǅ����    ������������������k�	�������������������������   3�tǅ����   �
ǅ����    ������������������ u!h��j ha  h�uj�o�������u̃����� uF腯���    j ha  h�uht�h��褦����ǅ��������M��0���������  ��������������������  �������$�0	�E�    �M��y���P������R�K���������   ������P�MQ������R�u  ���E��������U���U����������؉�|���u!h`tj h�  h�uj�m�������u̃�|��� uF胮���    j h�  h�uht�h`t袥����ǅ��������M��.���������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK��������h	�$�P	�E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�J������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�������Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ���������	�$�|	�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ���������	�$��	�U���0  u�E�   �E��M���  tUǅx���    �UR�ʟ����f������������Ph   ������Q�U�R�x�������x�����x��� t�E�   �&�EP�̧����f��t�����t����������E�   �������U��W  �EP蘧������p�����p��� t��p����y u�� �U��E�P�f������E��P�M���   t&��p����B�E���p�����+����E��E�   ��E�    ��p����B�E���p�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������h����MQ�Ŧ�����E��U���  te�}� u�� �E��E�   �M���d�����h�����h�������h�����t��d������t��d�������d����ɋ�d���+M����M��[�}� u	�� �U��E���l�����h�����h�������h�����t��l������t��l�������l����ɋ�l���+E��E��  �MQ��������`����O�������   3�tǅ����   �
ǅ����    ��������\�����\��� u!htj h�  h�uj�w�������u̃�\��� uF荨���    j h�  h�uht�ht謟����ǅ ��������M��8����� �����  ��  �U��� t��`���f������f����`�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h�sj�Ú�]  R�������E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���P�����T����M�袃��P�E�P�M�Q������R�E�P�M�Q��P���R��P��a�Ѓ��M���   t$�}� u�M��X���P�U�R��P��a�Ѓ���������gu*�U���   u�M��#���P�E�P��Q��a�Ѓ��U����-u�M���   �M��U����U��E�P�\������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�:�������@�����D����   �U���   t�EP��������@�����D����   �M��� tB�U���@t�EP�j���������@�����D�����MQ�N����������@�����D����=�U���@t�EP�(��������@�����D�����MQ������3҉�@�����D����E���@t@��D��� 7|	��@��� s,��@����ً�D����� �ډ�8�����<����E�   �E����@�����8�����D�����<����E�% �  u&�M���   u��8�����<����� ��8�����<����}� }	�E�   ��M�����M��}�   ~�E�   ��8����<���u�E�    �E��E��M̋Ũ��U̅���8����<���t{�E��RP��<���Q��8���R�b�����0��L����E��RP��<���P��8���Q�=�����8�����<�����L���9~��L����������L����E���L�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅4����M���u������R�EP��4���Qj �K	  ���U�R������P�MQ�U�R�E�P�|	  ���M���t$�U���u������P�MQ��4���Rj0� 	  ���}� ��   �}� ��   ǅ���    �E���0����M܉�,�����,�����,�������,�������   ��0���f�f������������Pj�� ���Q��(���R艣�����������0�������0�������� u	��(��� uǅ���������*�M�Q������R�EP��(���Q�� ���R�{  ���V�����E�P������Q�UR�E�P�M�Q�U  �������� |$�U���t������P�MQ��4���Rj ��  ���}� tj�E�P�\������E�    ����������� t������tǅ����    �
ǅ����   ���������������� u!h(�j h�  h�uj��}������u̃���� uC�����    j h�  h�uht�h(�������ǅ���������M�荡����������������������M��q����������M�3�萤����]ÍI ������/�|������	������!�*� �I 7������� ��C���]���Y�;� �V��MiD   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP蘑�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��j�h8�h5�d�    P���SVW�h1E�3�P�E�d�    �E������E�    j��q������u����C  j�v�����E�    �E�    �	�E���E�}�@��  �M�<� T �#  �U�� T�E��	�M؃�@�M؋U�� T   9E���   �M��Q����   �E؃x uaj
�u�����E�   �M؃y u.h�  �U؃�R�@b��u	�E�   ��E؋H���U؉J�E�    �   �j
�f�����Ã}� u+�E؃�P��b�M��Q��t�E؃�P��b�4����}� u-�M��A�U�������E����M�U�+� T��E��������}��t��   ��   h�   h��jj@j �{������E؃}� ��   �E�M؉� T��S�� ��S�	�E؃�@�E؋M�� T��   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃����� T�D�U�R�1p������u�E������������E������   �j������ËE܋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} ��   �E;�S��   �M���U������ T�<�um�=�/uB�M�M��}� t�}�t�}�t�(�URj��c��EPj��c��MQj��c�U���E������ T�U�3����\���� 	   �z���     �����]�����������������������������������������������������������̋�U��Q�} ��   �E;�S��   �M���U������ T�L����   �U���E������ T�<�th�=�/u<�U�U��}� t�}�t�}�t�"j j��c�j j��c�
j j��c�E���M������ T�����3����=���� 	   �oy���     �����]������������������������������������������������������������̋�U����}�u�y���     �˒��� 	   ����2  �} |�E;�Ss	�E�   ��E�    �M�M��}� u!h��j h;  h��j�Ko������u̃}� u<�x���     �Y���� 	   j h;  h��h��h���x���������   �E���M������ T�D
������؉E�u!hԮj h<  h��j�n������u̃}� u9�x���     �͑��� 	   j h<  h��h��hԮ�����������U���E������ T���]����������������������������������������������������������������������������������������������̋�U��j�hh�h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP�Db�E��}� u� bP�"l��������q  �}�u�M��@�M���}�u
�U���U�覒���E؃}��u�O����    �v���     ����#  �E�    �EP�M�Q蠔�����U���U�E����M؃����� T�E�D
�M����U؃����� T�L$�ဋU����E؃����� T�L$�E����M؃����� T�D
$$�M����U؃����� T�D$�E�   �E������   �K�}� u8�U����E؃����� T�T����E����M؃����� T�T�M�Q�di����Ã}� t�U؉U���E������EԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E���M����� T�M��E�   �U��z u_j
�l�����E�    �E��x u,h�  �M���Q�@b��u�E�    �U��B���M��A�E������   �j
��~����Ã}� t!�U���E������ T�TR��b�E�M�d�    Y_^[��]��������������������������������������������������������������������������̋�U��E���M������ T�D
P��b]������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    j�j�����E�    �EP�8�����f�E��E������   �j�}�����f�E�M�d�    Y_^[��]���������������������������������������������̋�U��Q�=)�u�e���=)�u���  �(j �E�Pj�MQ�)R��b��u���  �f�E��]��������������������������������̋�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M��ew���M���g������   t1�M���g��� ���   th��j jGhh�j�h������u̍M��g����z u*�} t�Ef��Uf�
�E�   �M������E��R  �M��gg��P�E�Q�:i��������   �M��Gg������   ~R�M��4g��� �M;��   |=3҃} ��R�EP�M��g������   R�EPj	�M���f����QR��a��uB�M���f��� �M;��   r�U�B��u"�[���� *   �E������M��'����E��   �M��f������   �U�M������E��k�a3��} ��P�MQj�URj	�M��hf��� �HQ��a��u����� *   �E������M�赊���E���E�   �M�衊���E���M�蔊����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�Ȇ����]�������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �E�    j�f�����E�    �E�   �	�E����E��M�;`S��   �U�@�<� t|�M��@���H��   t"�U�@��Q�#��������t	�U���U�}�|=�E��@���� R�Lbj�E��@��R�z�����E��@��    �Y����E������   �j�!y����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �} uj �  ���@�EP��t�����E�    �MQ�~�����E��E������   ��UR�|����ËE�M�d�    Y_^[��]������������������������������������������̋�U��} uj �n  ���@�EP�y�������t����+�M�Q�� @  t�EP�'q����P�hm��������3�]�����������������������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R�p����P�ڍ����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����������������������������������������������������̋�U��j�   ��]���������������̋�U��j�h�h5�d�    P���SVW�h1E�3�P�E�d�    �E�    �E�    j��b�����E�    �E�    �	�E����E��M�;`S��   �U�@�<� ��   �M��@���H��   ��   �U�@��Q�U�R�P������E�   �E��@���B%�   te�}u%�M��@��P�B{�������t	�M���M��:�} u4�U�@���Q��t!�E��@��R�{�������u�E������E�    �   ��E��@��R�E�P��x�����������E������   �j��t����Ã}u�E����E܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������̋�U����} uh(sj j?h�j��_������u̋M�M��U�R�m����P�G{������u3��  �tr���� 9E�u	�E�    ��^r����@9E�u	�E�   �3���   ��?����?�M��Q��  t3��   �E��<��? u\j[h��jh   �Z�����E�M��U���?�}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U����?�A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]��������������������������������������������������������������������������������������̋�U��Q�} t'�}t!h��j h�   h�j�"^������u̋M�M��} tG�U��B%   t:�M�Q�~�����U��B%�����M��A�U��B    �E��     �M��A    ��]��������������������������������������̋�U��j�h8�h5�d�    P���SVW�h1E�3�P�E�d�    �4p���� �E�3��} ���E؃}� uh(3j j4h��j�8]������u̃}� u+�Q����    j j4h��h��h(3�sw��������i�U�R��m�����E�    �E�P��������E܋MQ�UR�EP�M�Q�U���E��U�R�E�P�d|�����E������   ��M�Q�yu����ËE��M�d�    Y_^[��]�����������������������������������������������������������������������̋�U��EP�MQ�URh���ԅ����]����������������̋�U��EP�MQ�URh��褅����]����������������̋�U��EP�MQ�URhΝ�t�����]����������������̋�U��EPj �MQh���F�����]������������������̋�U��EPj �MQh��������]������������������̋�U��EPj �MQhΝ������]������������������̋�U���   �h3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���i���E�    ��}���E�3Ƀ} �������������� u!hLvj h  h�uj�Z������u̃����� uF�}���    j h  h�uhh�hLv�t����ǅ8��������M��I~����8����  3��} �������������� u!h(3j h  h�uj� Z������u̃����� uF�}���    j h  h�uhh�h(3�5t����ǅ4��������M���}����4����z  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���h  ������ �[  �������� |%��������x�������������� ����
ǅ ���    �� ���������������k�	�������������������������   3�tǅ���   �
ǅ���    ����������������� u!h��j ha  h�uj�X������u̃����� uF�{���    j ha  h�uhh�h����r����ǅ0��������M��S|����0����  �����������������*  ������$�\<�E�   ������Q�UR������P�Y  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ������������������ ����������wL��������<�$�|<�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�Aw�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP��v�����Ẽ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  ��������<�$��<�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  �������(=�$��<�M���0  u	�U��� �U��E�   �EP�u����f�������M��� tW���������   ������ƅ���� �M��oT��P�M��fT��� ���   Q������R������P�u������}�E�   �f������f�������������U��E�   �  �EP�t���������������� t�������y u�� �U��E�P�WX�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ�����������|����MQ�s�����E��U��� ��   �}� u�� �E��M��������E�    �	�U܃��U܋E�;�|���}L���������t?�M���R��P�������Q�T������t������������������������������d�}� u	�� �M��E�   �U���x�����|�����|�������|�����t��x������t��x�������x����ɋ�x���+U����U��  �EP�r������t����e������   3�tǅ���   �
ǅ���    �������p�����p��� u!htj h�  h�uj�DR������u̃�p��� uF�Zu���    j h�  h�uhh�ht�yl����ǅ,��������M��v����,����  ��  �M��� t��t���f������f����t�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h�sj�Ḿ�]  Q�L�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��oP��P�U�R�E�P������Q�U�R�E�P��h���Q��R��a�Ѓ��E�%�   t%�}� u�M��%P��P�M�Q��R��a�Ѓ���������gu)�M���   u�M���O��P�U�R��P��a�Ѓ��M����-u�E�   �E��M����M��U�R�*T�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�Y������X�����\����   �U���   t�EP��X������X�����\����   �M��� tB�U���@t�EP�2o��������X�����\�����MQ�o���������X�����\����=�U���@t�EP��n�������X�����\�����MQ��n����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R�'q����0��d����E��RP��T���P��P���Q�o����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �N  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��lK��P�M��cK������   R��H���P������Q�l������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�v  �������� |$�U���t������P�MQ��L���Rj ��  ���}� tj�E�P�-`�����E�    �s��������� t������tǅ ���    �
ǅ ���   �� �����<�����<��� u!h(�j h�  h�uj�J������u̃�<��� uC�m���    j h�  h�uhh�h(���d����ǅ(��������M��^n����(������������$����M��Bn����$����M�3��aq����]�h.�.�.8/�/�/�/1///�.*/3/ �I A0�00�0
1 ��4L1�2�6�1�4`1m6�3�6�6�26�6�9   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�n_�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����#  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tA�U�;U�u*�E�H�� ��Ƀ��U�� ��҃�;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �h3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T����N��ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �6b����|���3Ƀ} ����0�����0��� u!hLvj h  h�uj��>������u̃�0��� uI��a���    j h  h�uh��hLv�Y����ǅ,���������T����b����,����3  3��} ����,�����,��� u!h(3j h  h�uj�H>������u̃�,��� uI�^a���    j h  h�uh��h(3�}X����ǅ(���������T����b����(����3  ǅL���    �U������ǅ@���    ���@�������@�����@�����2  ��@���u������ u�2  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Mǅ��������ǅ��������ǅp�������ǅ���������Uf�f��D�����D����U���U���K/  ��L��� �>/  ��D����� |%��D�����x��D����������������
ǅ����    ��������H�����H���k�	��8����������8�����8�����  �U���%��  �������u\j
��t���Q�UR�B������~9��t������$u+��@��� uh@  j ������R�$h����ǅ����   �
ǅ����    �������)  j
��t���P�MQ�A��������������t������U��@��� ��   ������ |#��t������$u������d}ǅ����   �
ǅ����    ��������(�����(��� u!h8�j hQ  h�uj�c;������u̃�(��� uI�y^���    j hQ  h�uh��h8��U����ǅ$���������T����!_����$����40  ������;�x���~���������������x�����������������x����   ��8�����   3�tǅ����   �
ǅ����    ��������$�����$��� u!h��j h]  h�uj�{:������u̃�$��� uI�]���    j h]  h�uh��h���T����ǅ ���������T����9^���� ����L/  ��8����������������N,  �������$��{��@��� u	������t��@���u�������u�,  ǅ����   ��L���Q�UR��D���P�=  ����+  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �+  ��D����������������� ������������wj���������{�$��{���������������E���������������4���������������#�������ʀ   ����������������������	+  ��D�����*��  ������ u�UR�X�����������`  j
��t���P�MQ�4>��������������t������U��@��� ��  ������ |#��t������$u������d}ǅ|���   �
ǅ|���    ��|����� ����� ��� u!h(�j h�  h�uj��7������u̃� ��� uI�[���    j h�  h�uh��h(��-R����ǅ���������T����[���������,  ������;�x���~��������x������x�����x�����x�����x����������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R�bD��������؉����u!h��j h�  h�uj�6������u̃���� uI��Y���    j h�  h�uh��h����P����ǅ���������T����}Z��������+  �(  �+������������������������P�MV���������������� }���������������������ډ������������k�
��D����TЉ������2(  ǅd���    �#(  ��D�����*��  ������ u�MQ��U������d����`  j
��t���R�EP�N;��������p�����t������M��@��� ��  ��p��� |#��t������$u������d}ǅt���   �
ǅt���    ��t������������� u!h��j h�  h�uj�5������u̃���� uI�(X���    j h�  h�uh��h���GO����ǅ���������T�����X���������)  ��p���;�x���~��p�����p������x�����p�����p�����x�����p����������� uG��p�����Ǆ����   ��p�����f��D���f��������p������������������   ������Q��D���Rj��p�����������Q�|A��������؉����u!h �j h�  h�uj��3������u̃���� uI��V���    j h�  h�uh��h ��N����ǅ���������T����W��������(  ��%  �+��p���������������������R�gS������d�����d��� }
ǅd����������d���k�
��D����TЉ�d����_%  ��D�����l�����l�����I��l�����l���.�D  ��l�����|�$�|�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������d�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu������   �������ǅ8���    ������#�������� ���������������   ��������#  ��D�����h�����h�����A��h�����h���7�B!  ��h������|�$�H|��������0  u�������� ������ǅ����   ������ u�EP�BQ����f��<�����  ������ |������d}ǅd���   �
ǅd���    ��d������������� u!h��j hv  h�uj��0������u̃���� uI��S���    j hv  h�uh��h���K����ǅ���������T����T��������%  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�]=��������؉����u!hx�j hz  h�uj�/������u̃���� uI��R���    j hz  h�uh��hx���I����ǅ���������T����xS��������$  �  �,���������������� ����� ���Q�HO����f��<����������� t_��<���%�   ������ƅ���� ��T����.��P��T����.������   R������P��P���Q�O������}
ǅl���   �f��<���f��P�����P���������ǅ����   �^  ������ u�MQ�N������������  ������ |������d}ǅ`���   �
ǅ`���    ��`��������������� u!h��j h�  h�uj�$.������u̃����� uI�:Q���    j h�  h�uh��h���YH����ǅ���������T�����Q���������"  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�:��������؉�����u!h��j h�  h�uj�-������u̃����� uI�(P���    j h�  h�uh��h���GG����ǅ ���������T�����P���� �����!  �w  �+��������������������������R�L���������������� t�������x u#�� ������������R�h0�����������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q��������������������  ��������0  u�������� ��������d����uǅ\���������d�����\�����\��������������� u�EP�K������������  ������ |������d}ǅX���   �
ǅX���    ��X��������������� u!h��j h6  h�uj�%+������u̃����� uI�;N���    j h6  h�uh��h���ZE����ǅ����������T�����N����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�7��������؉�����u!h��j h:  h�uj�*������u̃����� uI�)M���    j h:  h�uh��h���HD����ǅ����������T�����M����������  �x  �+��������������������������Q�I������������������ ��   ������ u�� ������������������ǅ����    ���������������������;�����}O���������tB��T����(��P�������Q�}*������t������������������������������v������ u�� ������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������'  ������ u�EP�bH������������  ������ |������d}ǅT���   �
ǅT���    ��T��������������� u!h��j h�  h�uj��'������u̃����� uI�K���    j h�  h�uh��h���"B����ǅ����������T����K���������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�~4��������؉�����u!h��j h�  h�uj��&������u̃����� uI��I���    j h�  h�uh��h���A����ǅ����������T����J���������  �@  �+��������������������������Q�iF������������8������   3�tǅP���   �
ǅP���    ��P��������������� u!htj h�  h�uj��%������u̃����� uI�I���    j h�  h�uh��ht�/@����ǅ����������T����I����������  �_  �������� t������f��L���f����������L����ǅl���   �%  ǅh���   ��D����� f��D�����������@��������������  ��@��� ��  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u!h��j h�  h�uj��$������u̃����� uI��G���    j h�  h�uh��h����>����ǅ����������T����H���������  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R�e1��������؉�����u!h0�j h�  h�uj��#������u̃����� uI��F���    j h�  h�uh��h0���=����ǅ����������T����G���������  �'  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��D�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Yh�  h�sj��d���]  P�J���������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�E���E�M�Q��A��������������  ������ |������d}ǅH���   �
ǅH���    ��H��������������� u!h��j h  h�uj�"������u̃����� uI�0E���    j h  h�uh��h���O<����ǅ����������T�����E����������  ��@���t!h��j h  h�uj�!������u̋����������������������������������������Q��A���������������T����� ��P��h���Q��d���R��D���P��P���Q������R������P��Q��a�Ѓ���������   t.��d��� u%��T���� ��P������P��Q��a�Ѓ���D�����gu2������%�   u%��T����F ��P������Q��R��a�Ѓ����������-u!��������   ��������������������������Q�j$�����������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ������%�   t&�0   f��������4�����Qf������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  �%  ������ u�EP� )������������������  ������ |������d}ǅD���   �
ǅD���    ��D��������������� u!h��j h�  h�uj�
������u̃����� uI� B���    j h�  h�uh��h���?9����ǅ����������T�����B����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�+��������؉�����u!hH�j h�  h�uj��������u̃����� uI�A���    j h�  h�uh��hH��-8����ǅ����������T����A����������  �]  �1��������������������������Q�'�����������������  ��������   �%  ������ u�EP��&������������������  ������ |������d}ǅ@���   �
ǅ@���    ��@��������������� u!h��j h�  h�uj��������u̃����� uI��?���    j h�  h�uh��h���7����ǅ����������T����@���������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�d)��������؉�|���u!h��j h�  h�uj��������u̃�|��� uI��>���    j h�  h�uh��h����5����ǅ����������T����?���������  �&  �1����������������x�����x���Q��$������������������  �������� �e  ��������@�)  ������ u�MQ�;��������������������  ������ |������d}ǅ<���   �
ǅ<���    ��<�����t�����t��� u!h��j h�  h�uj�������u̃�t��� uI�=���    j h�  h�uh��h����4����ǅ����������T����L>���������_  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�'��������؉�p���u!hx�j h�  h�uj�|������u̃�p��� uI�<���    j h�  h�uh��hx��3����ǅ����������T����:=���������M  ��  �3����������������l�����l���R�
9�������������������(  ������ u!�EP��8���������������������  ������ |������d}ǅ8���   �
ǅ8���    ��8�����h�����h��� u!h��j h�  h�uj�c������u̃�h��� uI�y;���    j h�  h�uh��h���2����ǅ����������T����!<���������4  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P��$��������؉�d���u!hx�j h�  h�uj�Q������u̃�d��� uI�g:���    j h�  h�uh��hx��1����ǅ����������T����;���������"  �  �5����������������`�����`���Q��6��������������������Z  ��������@�'  ������ u�EP�6�������������������  ������ |������d}ǅ4���   �
ǅ4���    ��4�����\�����\��� u!h��j h  h�uj�*������u̃�\��� uI�@9���    j h  h�uh��h���_0����ǅ����������T�����9����������
  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�"��������؉�X���u!hx�j h  h�uj�������u̃�X��� uI�.8���    j h  h�uh��hx��M/����ǅ����������T�����8����������	  �}  �2����������������T�����T���Q�4������������������$  ������ u�UR�4����3ɉ�������������  ������ |������d}ǅ0���   �
ǅ0���    ��0�����P�����P��� u!h��j h0  h�uj�������u̃�P��� uI�7���    j h0  h�uh��h���7.����ǅ����������T�����7����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q� ��������؉�L���u!hx�j h4  h�uj��������u̃�L��� uI�6���    j h4  h�uh��hx��%-����ǅ����������T����6����������  �U  �3����������������H�����H���R�~2����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ��������������d��� }ǅd���   �%�����������������d���   ~
ǅd���   �����������u
ǅ����    ��O�����������d�����d�������d������������������   �������RP������P������Q�4����0�������������RP������R������P�p2��������������������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�k  ��l��� �:  ��������@tj��������   t�-   f������ǅ����   �D��������t�+   f������ǅ����   �!��������t�    f������ǅ����   ������+�����+�������D�����������u��L���Q�UR��D���Pj ��  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��D���Qj0�  �������� ��   ������ ��   ��������@�����������<�����<�����<�������<�������   ��T����F��P��T����:��� ���   Q��@���R��<���P�k/������8�����8��� ǅL��������2��L���Q�UR��<���P�E  ����@����8�����@����`����(��|���R��L���P�MQ������R������P��  ����L��� |'��������t��L���R�EP��D���Qj �T  �������� tj������R��"����ǅ����    ������8��� t��8���tǅ,���    �
ǅ,���   ��,�����4�����4��� u!h(�j h�  h�uj�_������u̃�4��� uI�u0���    j h�  h�uh��h(��'����ǅ����������T����1���������0  �������  ��@��� ��  ǅ����    ���������������������;�x�����  ����������������(�����(�������(�����(�����   ��(����$��|���������E�������MQ�t,�����_  ���������E�������MQ�P,�����;  ���������E�������MQ������  ���������E�������MQ�������   ���������E�������MQ��+������   ���������E�������MQ�s�����������������   3�tǅ$���   �
ǅ$���    ��$�����0�����0��� u!h��j h.	  h�uj�S������u̃�0��� uF�i.���    j h.	  h�uh��h���%����ǅ����������T����/���������'�����#�����L�����������T�����.���������M�3��2����]Ë��L�L&M�M�P�PdS�T�M�MpM_M�M�M �I �S�T�S�T�T �aU�Zgf�W7a0U0f^�f]f�ZNfsfAv   	
�y"zFzjz�z�z�z�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U��j�hX�h5�d�    P���SVW�h1E�3�P�E�d�    3��} ���E܃}� uh,�j j3h��j��������u̃}� u-����    j j3h��h��h,��>�������  �M�U�U�E�P�
�����E�    �M�Q�UR�����f�E��E������   ��E�P�_�����f�E��M�d�    Y_^[��]����������������������������������������������������������������������������̋�U���8�h3ŉE�V�E�H��@�d  �UR���������t@�EP��������t/�MQ����������UR���������� T�E���E���E�H$�����у�tj�EP�e�������t@�MQ�T�������t/�UR�C���������EP�2��������� T�E���E���M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ�"�����  �(  �UR��������t@�EP��������t/�MQ�q���������UR�`��������� T�E���E���E��H��   ��   �URj�E�P�M�Q��������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP� ����^�M�3��m����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ� ����]��������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���������������������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   �P��}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q��a_^��]� ���������������������̋�U��Q�M��E�� |��M��A    �U��B �E���]����������������������̋�U��Q�M��M������E��t�M�Q�f������E���]� �����������������̋�U��Q�M��E�� |��M��A    �U��B �E�Q�M��M����E���]� ���������������������̋�U��Q�M��E�� |��M��U��A�M��A �E���]� ������������������̋�U��Q�M��E�� |��M��A    �U��B �EP�M��y����E���]� �����������������������̋�U��Q�M��E�;Et0�M������M�Q��t�E�HQ�M��k�����U��E�H�J�E���]� ���������������������̋�U��Q�M��E�� |��M��z����]������������������̋�U����M��E��x t�M��Q�U���E����E���]�������������������̋�U����M��} tK�EP����������E��M�Q�������U��B�E��x t�MQ�U�R�E��HQ������U��B��]� �����������������������������̋�U��Q�M��E��H��t�U��BP�-�����M��A    �U��B ��]������������������������̋�U��Q�M��EP�M�����M�����E���]� ��������̋�U��Q�M��M��+����E��t�M�Q�v������E���]� �����������������̋�U��Q�M��EP�M��H���M�����E���]� ��������̋�U��Q�M��E�� ���M������]������������������̋�U��Q�M��EP�M��L���M�����E���]� ��������̋�U��Q�M��M������E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M��x���M�����E���]� ��������̋�U��Q�M��E�� ���M������]������������������̋�U��Q�M��EP�M������M�����E���]� ��������̋�U��Q�M��M������E��t�M�Q��������E���]� �����������������̋�U��Q�M��EP�M�������M�����E���]� ��������̋�U��Q�M��E�� ���M�� ����]������������������̋�U���8�EP�M�����3Ƀ} ���M�}� uh��j j4h��j�Q�������u̃}� u=�j���    j j4h��h��h��������E�����M�����E��  3��} ���E��}� uhL�j j5h��j���������u̃}� u=�����    j j5h��h��hL�������E�����M�����E��   �M��!�����z u"�EP�MQ�Z������EԍM��u���E��x�b�U��E̍M������P�M�Q��������E��U���U�E��MȍM�����P�U�R�������E��E���E�}� t�M�;M�t��U�+U��UЍM������EЋ�]����������������������������������������������������������������������������������������������������������̋�U����E��M��U��E���E��A|�}�Z	�M��� �M��U��E��M��U���U��A|�}�Z	�E��� �E��}� t�M�;M�t��E�+E���]������������������������������̋�U����=�? ��   3��} ���E��}� uh��j jbh��j��������u̃}� u0�����    j jbh��hh�h�������������   3҃} �U��}� uhL�j jch��j�J�������u̃}� u-�c���    j jch��hh�hL�����������&�MQ�UR���������j �EP�MQ��������]������������������������������������������������������������������������̋�U���@�} �!  �EP�M�����3Ƀ} ���M�}� uh��j j;h��j�W�������u̃}� u=�p���    j j;h��h��h��������E�����M��!���E��  3��} ���E��}� uhL�j j<h��j���������u̃}� u=�����    j j<h��h��hL�������E�����M�����E��1  ����;U����E�uh��j j=h��j�q�������u̃}� u=����    j j=h��h��h��������E�����M��;���E��   �M�������z u)�EP�MQ�UR��������E̍M�����E��   �m�E��MčM��r���P�U�R�o������E��E���E�M��U��M��H���P�E�P�E������E��M���M�U���Ut�}� t�E�;E�t��M�+M��MȍM��|���E��3���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����=�? �Y  3��} ���E��}� u!h��j h�   h��j��������u̃}� u3�
���    j h�   h��h@�h�������������  3҃} �U��}� u!hL�j h�   h��j�!�������u̃}� u3�:
���    j h�   h��h@�hL��Y���������   ����;M҃��U�u!h��j h�   h��j��������u̃}� u0��	���    j h�   h��h@�h���� ���������.�MQ�UR�EP�(�������j �MQ�UR�EP�e�������]��������������������������������������������������������������������������������������������������������̋�U��j j jj jh   @hX��c�)]����������̋�U��=)�t�=)�t�)P�c]�����������̋�U��j�hx�h5�d�    P���SVW�h1E�3�P�E�d�    �E�����3��} ���E��}� uhLvj j.h��j��������u̃}� u+�5���    j j.h��hl�hLv�W���������W�U�B��@t�M�A    �=�UR�������E�    �EP�e�����E��E������   ��MQ�o�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U����E�����3��} ���E�}� uh,�j jYh��j���������u̃}� u.����    j jYh��h��h,��1���������   �U�U��E��H��   ta�U�R������E��E�P�������M�Q�_�����P�������}	�E������$�U��z tj�E��HQ�}������U��B    �E��@    �E���]�����������������������������������������������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �}�u����� 	   ����  �} |�E;�Ss	�E�   ��E�    �M؉M��}� uh��j j,hp�j�_�������u̃}� u.�x��� 	   j j,hp�hX�h������������;  �E���M������ T�D
������؉E�uh�j j-hp�j���������u̃}� u.����� 	   j j-hp�hX�h������������   �UR��������E�    �E���M������ T�D
��t;�MQ������P�c��u� b�E���E�    �}� u�>�����U��a��� 	   �E�����3�uh �j jEhp�j��������u��E������   ��UR�P�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�   ��]�������������������̋�U���$�} t�E�M�3҃} �U�}� uh̼j j^h��j���������u̃}� u-�����    j j^h��hp�h̼������3��'  �} t�}|�}$~	�E�    ��E�   �M��M�}� uh�j j_h��j�`�������u̃}� u-�y���    j j_h��hp�h�������3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q���������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R�������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q�i������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q������E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4������ "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�X�����]�������������������̋�U��j�EP�MQ�UR�(�����]�������������������̋�U��j�EP�MQ�UR�������]�������������������̋�U��� �} uh(sj jdh�rj���������u̋M�M��U�R�������E��E��H��   u&������ 	   �U��B�� �M��A���  �c  �/�U��B��@t$����� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6������ 9E�t�~�����@9E�u�M�Q�-�������u�U�R�������E��H��  �  �U��E��
+Hy!hrj h�   h�rj�T�������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�&�����E��s�}��t!�}��t�M����U������ T�U���E���E��H�� t9jj j �U�R�7������E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q�r�����E�U�;U�t�E��H�� �U��J���  ��E%��  ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̋�U��j�h��h5�d�    P���SVW�h1E�3�P�E�d�    �}�u�����     ������ 	   ����  �} |�E;�Ss	�E�   ��E�    �M؉M��}� uh��j j.h�j�T�������u̃}� u9�����     �b���� 	   j j.h�h��h������������  �E���M������ T�D
������؉E�uhԮj j/h�j���������u̃}� u9�$����     ������ 	   j j/h�h��hԮ�����������   �UR��������E�    �E���M������ T�D
��t�MQ�g������E��4�j���� 	   �E�����3�uh �j j9h�j��������u��E������   ��MQ�Y�����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QV�EP�d��������t]�}u� T���   ��u�}u(� T�HD��tj�)�������j������;�t�UR������P�c��t	�E�    �	� b�E��EP�s������M���U������ T�D �}� t�M�Q�O���������3�^��]����������������������������������������������������̋�U��} uh��j j.h��j�,�������u̋M�Q��   tK�E�H��t@j�U�BP�(������M�Q�������E�P�M�    �U�B    �E�@    ]��������������������������������������������̋�U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%�a�%�a�%�a�%�a�%�a�%�a�%�a�%�a�%�a�%�a�% b�%b�%b�%b�%b�%b�%b�%b�% b�%$b�%(b�%,b�%0b�%4b�%8b�%<b�%@b�%Db�%Hb�%Lb�%Pb�%Tb�%Xb�%\b�%`b�%db�%hb�%lb�%pb�%tb�%xb�%|b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�%�b�% c�%c�%c�%c�%c�%c�%c�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̡d?����d?ËT$�B�J�3���������O�������������������������̍M��B����T$�B�J�3��`���������������������̍M������T$�B�J�3��0����(������������������̍M�������T$�B�J�3�� ����������������������̍M������T$�B�J�3������������������������̋T$�B�J�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫹄*葶��h ��������_^[���   ;��������]������������������������U����   SVW��@����0   ������j �`/跿��_^[���   ;�������]������������������̋�U��Q3��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫹄*�c���_^[���   ;��$�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                         0�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            7������Y�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��x�                                                                                                                                                                                                                                                                    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��P          �� �d
 IDM_NEU     SDK Test    IDS_EDITOR_PLUGINS      PLUGIN_CMD_1000472      M_EDITOR    C4DSDK - Edit Image Hook:       -plugincrash    -SDK executed:-)       -SDK    -SDK is here :-)       -help   --help  ����5�����a�:�ǆԃF�        MY BUTTON   MySecondGroup   &i  &   MyGroup     MyTextGroup     Hello       �������        ������              �?                    Custom GUI Button Was Pressed       Fouth Option Selected       Third Option Selected       Second Option Selected      First Option Selected       CHKBox was Toggled      icon error      Button Was Pressed          .   C++ RES Based Dialog        icon.tif    c:\program files\maxon\cinema 4d r12\plugins\resbaseddialog_c++\source\myresdialog.cpp                  C++ Dialog using external resources         res myicon.png      �� �h��G�L���x�        ����Q���L�\��x�        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp                 #   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp                %s      c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h                ��R�������Ռa�:�ǆT�             �f@        -DT�!	@              Y@             @�@    ����������Ռa�:�ǆ��        $���ɱ2�g�`�T�>�����Z�J�            c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gui.cpp              |���������Ռa�:�ǆ`�        ~   ��E�������Ռa�:�ǆ��L�֩f�q�V���9�~���<���ر                    Progress Thread     0%  %   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_memory.cpp               c:\program files\maxon\cinema 4d r12\resource\_api\c4d_string.cpp               no baselist      B   KB  MB           �@     GB c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp               8��    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp                      �?          4&�k�          4&�kC        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basetime.cpp                      �Ngm��C           ����A        ����MbP?    P�������    ���    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp                  �=�    ���    ��8�    �>�    c:\program files\maxon\cinema 4d r12\resource\_api\ge_sort.cpp              d��     �    f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c            f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c                   �?      �?3      3            �      0C       �       ��                                                          fmod         �fp	�o	fp	�o	fp	�o	fp	�o	�o	'p	�o	fp	fp	�o	fp	                Unknown Runtime Check Error
       Stack memory around _alloca was corrupted
         A local variable was used before it was initialized
           Stack memory was corrupted
            A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                �	@���                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                  Run-Time Check Failure #%d - %s         Unknown Module Name     Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s                   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                           Stack corrupted near unknown variable               Stack area around _alloca memory reserved by this function is corrupted
                %s%s%s%s    >   
   %s%s%p%s%ld%s%d%s           Stack area around _alloca memory reserved by this function is corrupted                 
Address: 0x    
Size:      
Allocation number within this function:            
Data: <    wsprintfA   u s e r 3 2 . d l l         %.2X    A variable is being used without being initialized.             Stack around _alloca corrupted          Local variable used before initialization           Stack memory corruption     Cast to smaller type causing loss of data           Stack pointer corruption        ���l    f:\dd\vctools\crt_bld\self_x86\crt\prebuild\misc\i386\chkesp.c                  The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p                             p N o d e - > _ N e x t   ! =   N U L L                 s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                 _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                       _ s e t d e f a u l t p r e c i s i o n                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c                         s i z e I n B y t e s   >   0           _ c f t o e _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c                         b u f   ! =   N U L L       e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                           _ c f t o e 2 _ l           s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o a _ l         _ c f t o f _ l         _ c f t o f 2 _ l       _ c f t o g _ l         f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c           FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    K E R N E L 3 2 . D L L         Client  Ignore  CRT Normal  Free    4,(     Error: memory allocation: bad memory block type.
           Invalid allocation size: %Iu bytes.
        Client hook allocation failure.
        Client hook allocation failure at file %hs line %d.
                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c                         _ C r t C h e c k M e m o r y ( )           _ p F i r s t B l o c k   = =   p O l d B l o c k               _ p L a s t B l o c k   = =   p O l d B l o c k             f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       Error: possible heap corruption at or near 0x%p                 p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Client hook re-allocation failure.
         Client hook re-allocation failure at file %hs line %d.
             _ e x p a n d _ d b g       p U s e r D a t a   ! =   N U L L           _ p F i r s t B l o c k   = =   p H e a d           _ p L a s t B l o c k   = =   p H e a d             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                                 HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()                _ m s i z e _ d b g         %hs located at 0x%p is %Iu bytes long.
             %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
                   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 DAMAGED     _heapchk fails with unknown return value!
          _heapchk fails with _HEAPBADPTR.
       _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADBEGIN.
         _ C r t S e t D b g F l a g             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t D o F o r A l l C l i e n t O b j e c t s               p f n   ! =   N U L L       Bad memory block found at 0x%p.
        Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              _ C r t M e m C h e c k p o i n t           s t a t e   ! =   N U L L           n e w S t a t e   ! =   N U L L         o l d S t a t e   ! =   N U L L         _ C r t M e m D i f f e r e n c e           Object dump complete.
      crt block at 0x%p, subtype %x, %Iu bytes long.
             normal block at 0x%p, %Iu bytes long.
          client block at 0x%p, subtype %x, %Iu bytes long.
              {%ld}   %hs(%d) :       #File Error#(%d) :      Dumping objects ->
      Data: <%s> %s
     ( * _ e r r n o ( ) )       _ p r i n t M e m B l o c k D a t a             Detected memory leaks!
     Total allocations: %Id bytes.
          Largest number used: %Id bytes.
        %Id bytes in %Id %hs Blocks.
       _ C r t M e m D u m p S t a t i s t i c s           o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g               Damage before 0x%p which was allocated by aligned routine
                  The block at 0x%p was not allocated by _aligned routines, use realloc()                 The block at 0x%p was not allocated by _aligned routines, use free()                _ a l i g n e d _ m s i z e _ d b g             m e m b l o c k   ! =   N U L L         CorExitProcess      m s c o r e e . d l l       _ w p g m p t r   ! =   N U L L         _ g e t _ w p g m p t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 d a t . c                         p V a l u e   ! =   N U L L         _ p g m p t r   ! =   N U L L           _ g e t _ p g m p t r       f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c             s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               _ s e t e n v p             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c            f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c            f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c          f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h e a p i n i t . c                       _ c r t h e a p           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                                      �1�1        ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                 _ v s n p r i n t f _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c                       ( f o r m a t   ! =   N U L L )               �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��                    tan cos sin modf    floor   ceil    atan    exp10   acos    asin    pow exp log10   log _nextafter      _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    �������             ��      �@      �                               ���5�h!����?      �?          r u n t i m e   e r r o r            
     T L O S S   e r r o r  
           S I N G   e r r o r  
         D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                            �>   P>	   �=
   �=   =   �<   X<   �;   p;   ;   �:   :   �9   h9   x8    �7!   �5x   �5y   d5z   @5�   85�   5                                        M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             
 
     w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                               . . .       w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           < p r o g r a m   n a m e   u n k n o w n >             w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                             R u n t i m e   E r r o r ! 
 
 P r o g r a m :                     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     _ N M S G _ W R I T E           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c                         s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         _ _ g e t l o c a l e i n f o               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t h e l p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\inithelp.c           M S P D B 1 0 0 . D L L     M S V C R 1 0 0 D . d l l               r   PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y                 S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S                       RegCloseKey     RegQueryValueExW    RegOpenKeyExW   A D V A P I 3 2 . D L L         D L L       M S P D B 1 0 0         ... Assertion Failed    Error   Warning     �G�G�G    f:\dd\vctools\crt_bld\self_x86\crt\src\dbgrpt.c             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       p f n N e w H o o k   ! =   N U L L             _ C r t S e t R e p o r t H o o k 2                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c                           m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           Microsoft Visual C++ Debug Library          _CrtDbgReport: String too long or IO Error          s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                     Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)                    
Module:    
File:      
Line:      

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.                              m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                 <program name unknown>      s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         _ _ c r t M e s s a g e W i n d o w A           A s s e r t i o n   F a i l e d         E r r o r       W a r n i n g       4N$N�M    _ C r t S e t R e p o r t H o o k W 2           M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y                     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )                                     
 M o d u l e :         
 F i l e :         
 L i n e :         E x p r e s s i o n :               
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                     w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       _ _ c r t M e s s a g e W i n d o w W           f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c          ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               B u f f e r   i s   t o o   s m a l l           ( ( ( _ S r c ) ) )   ! =   N U L L             s t r c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                      Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete      new    __unaligned     __restrict      __ptr64     __eabi  __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(        8[,[ [[[�Z�Z�Z�Z�Z�Z��Z�Z�Z�Z�Z�Z�Z�Z�ZxZtZpZlZhZdZ`Z��\ZXZ�TZPZLZHZDZ@Z\<Z8Z4Z0Z,Z(Z$Z ZZZZZZZ�Y�Y�Y�Y�Y�Y�YtYPY,YY�X�X�XpXHXX�W�W�W�W�W�W�W�WpWPW,W�V�V�VlVLV$V�U�U�UlU�TU0UU�T�T                                                                                CV:     ::  '   `   generic-type-   template-parameter-     ''  `anonymous namespace'       `non-type-template-parameter        `template-parameter     void    NULL    extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{    }'  }'  )   void    std::nullptr_t      volatile    ,<ellipsis>     ,...    <ellipsis>       throw(      volatile   const   signed      unsigned    UNKNOWN     __w64   wchar_t     <unknown>   __int128    __int64     __int32     __int16     __int8  bool    double  long    float   long    int short   char    enum    cointerface     coclass     class   struct      union   `unknown ecsu'      int     short   char    const   volatile    cli::pin_ptr<   cli::array<     )[  {flat}  s   {for    ���    ����}�    �����    �����    ���!�     ??     ��e�d�    _ c o n t r o l f p _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c                           ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c                       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )                                                                                         H H : m m : s s         d d d d ,   M M M M   d d ,   y y y y           M M / d d / y y         P M     A M     D e c e m b e r         N o v e m b e r         O c t o b e r       S e p t e m b e r       A u g u s t     J u l y     J u n e     A p r i l       M a r c h       F e b r u a r y         J a n u a r y       D e c       N o v       O c t       S e p       A u g       J u l       J u n       M a y       A p r       M a r       F e b       J a n       S a t u r d a y         F r i d a y     T h u r s d a y         W e d n e s d a y       T u e s d a y       M o n d a y     S u n d a y     S a t       F r i       T h u       W e d       T u e       M o n       S u n       HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun p f l t   ! =   N U L L             s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           _ f p t o s t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c                       _ g e t _ e r r n o             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d o s m a p . c                       _ g e t _ d o s e r r n o           s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                     _ f l t o u t 2             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c                         _ s e t _ o u t p u t _ f o r m a t             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t f o r m a t . c                               ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h a n d l e r . c p p                         p n h   = =   0         _ e x p a n d _ b a s e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c                       p B l o c k   ! =   N U L L         ( s t r i n g   ! =   N U L L )         s p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c                         ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6             s i g n a l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c                       ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f:\dd\vctools\crt_bld\self_x86\crt\src\winsig.c             r a i s e       SystemFunction036           ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       r a n d _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r a n d _ s . c                       _ R a n d o m V a l u e   ! =   N U L L             ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c                         s t r   ! =   N U L L       ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c             ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 ( c h   ! =   _ T ( ' \ 0 ' ) )         (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       _ o u t p u t _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c                       ( s t r e a m   ! =   N U L L )         _ s e t _ e r r o r _ m o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c                         ( " I n v a l i d   e r r o r _ m o d e " ,   0 )               GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L             ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               w c s c a t _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                     w c s n c p y _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l                         w c s c p y _ s         s t r n c p y _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h                           ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                   _ w m a k e p a t h _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t m a k e p a t h _ s . i n l                         ( L " I n v a l i d   p a r a m e t e r " ,   0 )               _ w s p l i t p a t h _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t s p l i t p a t h _ s . i n l                           ( ( ( _ P a t h ) ) )   ! =   N U L L           f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t M o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c                         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   _ C r t S e t R e p o r t F i l e               _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       %s(%d) : %s         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed!       Assertion failed:           s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   , Line      <file unknown>      Second Chance Assertion Failed: File            _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t A           w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               _CrtDbgReport: String too long or Invalid characters in String                  s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       % s ( % d )   :   % s       w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                 w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d !           A s s e r t i o n   f a i l e d :                   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 
   ,   L i n e         < f i l e   u n k n o w n >             S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t W           GetUserObjectInformationA       MessageBoxA     s i z e I n B y t e s   > =   c o u n t             s r c   ! =   N U L L       m e m c p y _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c                       d s t   ! =   N U L L       _ s w p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s w p r i n t f . c                            _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                         _ s e t _ c o n t r o l f p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                             LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL  8�    �(�<|��<%��<����<���<��                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         _ c o n f i g t h r e a d l o c a l e           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t l o c a l . c                       ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                       f:\dd\vctools\crt_bld\self_x86\crt\src\setlocal.c           s e t l o c a l e       L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     s t r n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ s e t l o c a l e _ n o l o c k           ;   =;  s t r c p y _ s ( p c h   +   s i z e o f ( i n t ) ,   c c h   -   s i z e o f ( i n t ) ,   l c t e m p )                         _ s e t l o c a l e _ s e t _ c a t             s t r c a t _ s ( p c h ,   c c h ,   " ; " )               _ s e t l o c a l e _ g e t _ a l l             s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   s t r n c p y _ s ( c a c h e i n ,   c a c h e i n S i z e ,   s o u r c e ,   c h a r a c t e r s I n S o u r c e   +   1 )                               C   s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   " C " )                 _ e x p a n d l o c a l e           s t r c a t _ s ( o u t s t r ,   s i z e I n B y t e s ,   (   * ( c h a r   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                           _ s t r c a t s             s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                               s t r n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   l o c a l e ,   l e n )                                             s t r n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                           _., s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & l o c a l e [ 1 ] ,   1 6 - 1 )                                             _ _ l c _ s t r t o l c         _       s t r c p y _ s ( l o c a l e ,   s i z e I n B y t e s ,   ( c h a r   * ) n a m e s - > s z L a n g u a g e )                         _ _ l c _ l c t o s t r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t t i m e . c                       p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                   f:\dd\vctools\crt_bld\self_x86\crt\src\inittime.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t n u m . c                         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initnum.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t m o n . c                         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initmon.c                                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                            _ _ s t r g t o l d 1 2 _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l                             _ L o c a l e   ! =   N U L L           1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 $ I 1 0 _ O U T P U T       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c                             _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r           _ v s n p r i n t f _ h e l p e r           ( " B u f f e r   t o o   s m a l l " ,   0 )               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   _ v s p r i n t f _ s _ l           f o r m a t   ! =   N U L L         _ v s n p r i n t f _ s _ l         ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   ( _ o s f i l e ( f h )   &   F O P E N )           _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c                       ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c                     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )               ( ( c n t   &   1 )   = =   0 )         _ w r i t e _ n o l o c k           ( b u f   ! =   N U L L )           f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c                         _ i s a t t y           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c          _ f i l e n o       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c                       p r i n t f         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p r i n t f . c                       _ w c t o m b _ s _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c                       s i z e I n B y t e s   < =   I N T _ M A X             _ m b s t o w c s _ l _ h e l p e r                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c                       s   ! =   N U L L       r e t s i z e   < =   s i z e I n W o r d s             b u f f e r S i z e   < =   I N T _ M A X           _ m b s t o w c s _ s _ l           ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                               s t r c a t _ s         l e n g t h   <   s i z e I n T C h a r s           2   < =   r a d i x   & &   r a d i x   < =   3 6               s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   s i z e I n T C h a r s   >   0         x t o a _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c                       x 6 4 t o a _ s         _ w c s t o m b s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c                       p w c s   ! =   N U L L         s i z e I n B y t e s   >   r e t s i z e           _ w c s t o m b s _ s _ l           ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               _ v s w p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c                       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s w p r i n t f _ s _ l         _ v s n w p r i n t f _ s _ l           x t o w _ s     x 6 4 t o w _ s         _ w o u t p u t _ l         _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r                 i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                   s t r t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o l . c                       n p t r   ! =   N U L L         s t r t o x q       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o q . c                       Ǥbad exception   ��[�ѩ    p l o c i - > c t y p e 1 _ r e f c o u n t   >   0             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t c t y p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\initctyp.c           united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american    T�ENU @�ENU ,�ENU �ENA �NLB �ENC  �ZHH ��ZHI ��CHS ��ZHH ��CHS ��ZHI ��CHT ��NLB p�ENU `�ENA L�ENL <�ENC $�ENB �ENI  �ENJ ��ENZ ��ENS ��ENT ��ENG ��ENU ��ENU p�FRB \�FRC D�FRL 4�FRS  �DEA �DEC ��DEL ��DES ��ENI ��ITS ��NOR ��NOR ��NON l�PTB T�ESS @�ESB 0�ESL �ESO �ESC ��ESD ��ESF ��ESE ��ESG ��ESH x�ESM d�ESN L�ESI 8�ESA $�ESZ �ESR ��ESU �ESY пESV ��SVF ��DES ��ENG ��ENU ��ENU                                                                                                         ��USA ��GBR ��CHN ��CZE t�GBR d�GBR X�NLD L�HKG <�NZL 8�NZL ,�CHN  �CHN �PRI �SVK ��ZAF �KOR ؾZAF ȾKOR ��TTO ��GBR ��GBR ��USA ��USA                                     6-    Norwegian-Nynorsk           s t r c p y _ s ( l p O u t S t r - > s z L a n g u a g e ,   ( s i z e o f ( l p O u t S t r - > s z L a n g u a g e )   /   s i z e o f ( l p O u t S t r - > s z L a n g u a g e [ 0 ] ) ) ,   " N o r w e g i a n - N y n o r s k " )                                                   _ _ g e t _ q u a l i f i e d _ l o c a l e                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t q l o c . c                         OCP ACP ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 _ o u t p u t _ p _ l           ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f:\dd\vctools\crt_bld\self_x86\crt\src\osfinfo.c            _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c                           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                             f:\dd\vctools\crt_bld\self_x86\crt\src\_sftbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ s f t b u f . c                         f l a g   = =   0   | |   f l a g   = =   1             v p r i n t f _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v p r i n t f . c                         _ w o u t p u t _ s _ l         _ w o u t p u t _ p _ l         f p u t w c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t w c . c                       ( s t r   ! =   N U L L )           csm�               �                X�m�ѩ    Unknown exception       p�?�ѩ    ����ѩ    (��ѩ    _ s t r i c m p _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r i c m p . c                         _ s t r i c m p         c o u n t   < =   I N T _ M A X         _ s t r n i c m p _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c m p . c                       _ s t r n i c m p       C O N O U T $       f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c                       _ f c l o s e _ n o l o c k         ( _ o s f i l e ( f i l e d e s )   &   F O P E N )             _ c o m m i t           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c                           ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         w c s t o x l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o l . c                       _ c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c                     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c                       s t r e a m   ! =   N U L L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             RSDS
���\��J�� ��(    C:\Program Files\MAXON\CINEMA 4D R12\plugins\ResBasedDialog_C++\obj\ResBasedDialog_C++_Win32_Debug.pdb                                                                                                                                                                                                                                                                                                       0�               D�    P�t�            ����    @   0�                ����    @   ��                   ��    t�                <��               ��    ���X�    <       ����    @   ��        \       ����    @   8�                   L�    �X�    |        ����    @   |�                   ��    X�                \8�                ��                ���               ��     �t�    �       ����    @   ��                    �<�               P�    X�    �        ����    @   <�                    ���               ��    ��t�    �       ����    @   ��                    ��               �    ���t�           ����    @   ��                    ||�                dh�               |�    ��    d        ����    @   h�                    ���               ��    ��    �        ����    @   ��                    ��               ,�    8�\�    �       ����    @   �        �        ����    @   ��                   ��    \�                ���                ���               ��    ��    �        ����    @   ��                    $�               8�    @�            ����    @   $�                    @|�               ��    ��    @        ����    @   |�                    �$��               ��    ���    �$       ����    @   ��        %        ����    @   <�                   P�    �                %<�                �(��               ��    ���    �(       ����    @   ��                    �(��               ��    ��    �(       ����    @   ��                    �(@�               T�    d���    �(       ����    @   @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ލލލލލލލލލލލލލލލލލލލލލލ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌڌ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����    ����    ����    '�    ����    ����    ����5�P�    ����    ����    ����    K�    ����    ����    ����D�J�    ����    ����    ������    ����    ����    ����    �    ����    ����    ����     �    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    4�    ����    ����    ����    "�����    y�        ����    ����    ����    h�����    ��        ����    ����    ����    |�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    q�    ����    ����    ����    ��    ����    ����    ����    F�    ����    ����    ����    U�    ����    ����    ����    � 	    ����    ����    ����    >	    ����    ����    ����    �	    ����    ����    ����    {	    ����    ����    ����    �	    ����    ����    ����    n#	    ����    ����    �����i	�i	    ����    ����    ����    �	    ����    ����    ����    ��	    ����    ����    ����    �	    ����    x���    ����    �	    ����    x���    ����    ӟ	    ���� �"�   ��                           ����    ����    ����    Qp
    ����    ����    ����    s
    ����@�"�   �                           ����    ����    ����    ��
    ����    ����    ����	�
#�
    ����    ����    �����
�
    ����    ����    �����
�
    ����    ����    ����    �
    ����    ����    ����    ��
    ����    ����    ����    ��
    ����p�"�    �                           ����    ����    ����    �        E        ����    |��    ����    �        Z        ����    ����    ����    �D    ����    ����    ����    �E����    F        ����    ����    ����    bJ����    �J        ����    ����    ����    GM        LL        M            ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ������"�   ��                           ����л"�    �                               ��    D�       T�t�        �$    ����       կ        %    ����       M�        ����    ����    ����    -c    �b
c        ����    ����    ����    �f    �e�e        ����    ����    �����j�j    ����    ����    �����l�l    ����    ����    ����sm~m    ����    ����    ����+u8u    ����    ����    �����u�u    ����    ����    ����lvyv    ����    ����    ����w%w    @           �x����    ����                  ��"�   ��   ��                       ����    ����    ����    �        s        ����    ����    ����    3    ����    ����    ����    �    ����    ����    ����    "    ����    ����    ����    �!    ����    ����    ����    �"    ����    ����    ����    �%        �%        ����    ����    ����    �)    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    |�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��P    b          X \ ` J� y   ResBasedDialog_C++.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   .?AVmyDialog@@          .?AVGeDialog@@      �       .?AVmyResDialog@@           .?AVCommandData@@           .?AVBaseData@@      8   Y  �  @      .?AVGeModalDialog@@             .?AVGeUserArea@@          u      .?AVSubDialog@@         .?AViCustomGui@@        c  �  �   �      �   �   �  �  Q      (   2       .?AVC4DThread@@         .?AVGeToolDynArray@@        -       .?AVGeToolDynArraySort@@            .?AVGeSortAndSearch@@           .?AVGeToolList2D@@          .?AVGeToolNode2D@@      �               .?AVtype_info@@     u�  s�      N�@���D                   '�'�'�'�'�'�'�'�'�'�        ��������       ����   ��������        �����
                                                                      ?     4   4    4   4   �4   �4!   �4   4    4   �3   �4   x4   �3   �3    �3   �3   �3   p4   �3   h4   `4   X4   P4   H4"   D4#   @4$   <4%   44&   $4                                                      �      ���������              �               �D        � 0                    �G�A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ����C   �h�h�h�h�h�h�h�h�h�h�h�h|hphlhhhdh`h\hXhThPhLhHhDh@h4h(h hh\hhh h�g�g�g�g�g�g�g�g�g	         �g�gtghg\gPgDg4g$gg�f�f�f�f�f�f�f�f|fpfdfXfLf@f4f(ff�e�e�e|f�e�e�e�e�epeXePeHe0e e�d                                                                                                                                                                   <            <            <            <            <                              @!        ���� �@                                            ��                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                         ��            TsDs    �&  ����         ������������                     �                ��.   .   8!�?�?�?�?�?�?�?�?�?<!�?�?�?�?�?�?�?@!                    ����       ���5      @   �  �   ����                         `C    `C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 .?AVbad_exception@std@@             .?AVexception@std@@                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                        .?AVbad_cast@std@@          .?AVbad_typeid@std@@            .?AV__non_rtti_object@std@@         ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (`         di �a                     �c �c �c �c �c �c �c d "d .d @d Pd \d jd xd �d �d �d �d �d �d �d 
e e (e :e Je re �e �e �e �e �e �e f f *f :f Pf jf ~f �f �f �f �f �f 
g g (g 4g Fg Vg dg |g �g �g �g �g �g �g �g �g �g h .h Dh Zh jh �h �h �h �h �h �h �h �h i $i 4i Bi Pi                                                                                                             �c �c �c �c �c �c �c d "d .d @d Pd \d jd xd �d �d �d �d �d �d �d 
e e (e :e Je re �e �e �e �e �e �e f f *f :f Pf jf ~f �f �f �f �f �f 
g g (g 4g Fg Vg dg |g �g �g �g �g �g �g �g �g �g h .h Dh Zh jh �h �h �h �h �h �h �h �h i $i 4i Bi Pi                                                                                                             �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer WideCharToMultiByte  IsDebuggerPresent gMultiByteToWideChar �RaiseException  MlstrlenA  EGetProcAddress  ?LoadLibraryW  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  GetLastError  �InterlockedDecrement  �GetCurrentThread  �HeapValidate  �IsBadReadPtr  ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter IsProcessorFeaturePresent GetModuleFileNameW  %WriteFile GetLocaleInfoW  �HeapFree  �HeapAlloc JGetProcessHeap  �VirtualQuery  bFreeLibrary � EnterCriticalSection  9LeaveCriticalSection   FatalAppExitA RtlUnwind hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage �HeapReAlloc �HeapSize  �HeapQueryInformation  -SetConsoleCtrlHandler �InterlockedExchange �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -LCMapStringW  iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  GetLocaleInfoA  IsValidLocale EnumSystemLocalesA  �GetUserDefaultLCID  �SetStdHandle  � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 � D   �5�5Q6�6�6�697�7Y8|8�8[9�9:�:�;<�<==�=�=�=|>�>�>?N?~?�? � L   0s1�1�1�123�3 4�4Q5�5\6n6D7V7,8>89&9:h:�: ;;;$;0;<;�=?>�>�?     P   0h0�23@3z3�3�34M4�4�45(545@5�67{7[8�8�9�9�9�9�9�9�9�:K;<�<=�=%>    D   0/011"1+1h1z1242@2L2X2�3`47�78�8�9/:�:�;<�<O>�>;?�?     X   @0�1�3�3�3R45�5<6T6�67c7x7888D8P8�8_9�9�9l:;,;8;D;�;�;|< =�=�=�=�=�>�>,?�?   0 `   40�0�0 11�1k2�3�3�3�3�3�45n6�6�6�6�6{7u8�8�8�8�8?9�9�9:�:�:3;U;�;<�<=�=>t>�>b?�?   @ L   �0"1;2�23�34�45�5�5�56o6�6o7�7o8�8F9�9/:�:.;�;<�<=�=>�>�>d?�? P D   K0�0+1�12{2�2[3�3�:�:�:O;t;�;�;'<�<= =�=�=�=�>�>�>S?x?�?   ` L   0�0�1�1l2�2K3�3;4�4-5�5�5�6&7�7�7h8�8^9�9�:;x;�;d<�<D=�=$>�>?�?   p L   0�0�0m1�1M2�2*3�3�4�4�4v5�5f6�6V7�798�8Z9�9�9�:�;&<�<$=�=>{>�>[?�? � P   ;0�01�1�1k2�2K3�3+4�45{5�5[6�6O7�7K8�8r9�9|:�:\;�;;<�<=�=>�>?{?�?   � L   [0�0;1�12�2�2w3�3_4�4g5�5T6�6;7�78�89�9�9d:�:b;�;z<�<_=�=?>�>7?�? � X   +0�0.1�1B2�2G3�3R4�4O5�5J6�6*7�78~8�8�8�8/9�9�9_:�::;�;<�<==�=v>�>U?�?�?�?�? � X   60�011�1?2�23�3�3r4�4Z5�56(646�6
7�7�7_8�869�9:T:x:�:�:F;�;j<�<m=�=M>�>-?�? � `   
0z0�0V1�1G2q2�2�2�2�273a3�3�3�3�3'4Q4t4�4�4�45�5�678�89�9:o:�:V;�;/<�<�<f=�=R>�>U? � \   0�01 1�1�1p2�2�34�4�4�56�697�7/8d8j8�8�8�8k9p9�9i:�:�;<<�<=(=>,>8>?4?@?�?   � T   0�0�0)1�12�23v3�3]4�4=5�56�6�6m7�7f8�8F9�9-:�:;z;�;V<�<=�=�=m>�>$?0?�? � D   0�0h4s4y45�5�5(6L6X6h7�78�89�90:�:t;�;�;�;�;o<=K=�=�>     8   !0�0`1�1�2K34�4;5N7t7�7&9L9X9�9	;0;<;<=<=H=�=  `   C0I0�0�0�0�1@2p2�2�203�3*5�5�5�5'7L7X7�7�8�8�8O9t9�9:,:8:�:$;0;�;�<�<�<�=�=�=>�>? ?,?   4   0�1�57�79�9�9�:B;Q;�;�;�;%=�=>>>+?�?   0 �   0(040�0j1�1�1�1Z2|2�2�2D3 4"4H4T4�4585D5�56(646�6�67$7�7`8�8�8�8P9r9�9�9@:b:�:�:0;R;x;�;<@<h<t<=0=X=d=�= >H>T>�>?8?D?�?   @ d   0(040�0�01$1�1p2�2�2�2`3�3�3�3N4p4�4�4?56@6L6X6d67�7�788�839�9C:�:^;�;~<�<�=1>�><?\?�? P @   �01�1W2�2�3�34$4�4^5�5�6:7�7�7�8 9�9@:�:f; <�<D=�=p>   ` P   �0�1 5 66666666 6�6084888<8@8D8H8L8P8x:X;p;<�<�<�<n=�=N>�>.?�?   p \   M01	1�12�23�3"4�415�566�6,8T8`8l8x8�8�8�8Q9�9V:�:F;�;F<�<n=�=�=�=>`>y>~>�>�>m?   � ,   0�0.1�12�263�3�4v567�7*8�8�;$=? � 0   B0h0t0�0�2h3�4F5�5�6'7L7X7�7Y8<=�=:>�>.? � 0   �5�5�5 666$606�7;9�9":�:@;�;�<1=�?�?�? � @   �0�0�0�1�1�1�2�2�2�3�3�3�4�4�4P6x6�6�7 8,8Q9x9�9 :>@>L> � 0   �05!6&6�6�6�78~8�89+:0:Y:�:�:3<X<d<R? � ,   �8&9�9
:z:�:�;�;�<=A=�=>�>�>\?�?�? � H   %0�01p1�102o2�2m3�3�3�3]4y4�4�4�4�5�5f6�6F7�708�829�9/:O;�<�<�< � X   {0�0�0�0�0�1�1�1�1W2m2r22�2T3�3�3F4l4�4w5�5�5J6�6�6!7{7�7�79O:�<=�=�={>�>k?�?   L   ;0�01�1�1h2�2�34�4�4k5�5_6�6k7�7K8�8;9�9K:�:/;�;/<�</=�=+>�>??�?  D   r0�0q1�1q2{3�3�3"6�78(8�8�9�9�9�:�:�:k;k<�<�<�=�=�=[>�>G?�?   4   61\1h1v2�2�2�3�3�3�455R8v<�<�<�=�=�=�>?? 0 D   f2�2?3�34�45?5�5�6.7�78�89�9:�:�;?<�<�<�<�<">�>?�?�?   @ L   k0�0[1�1?2�2�2�2�23+5�5+6�67�78�89):L:X:d:y;�;�;�;=<�<==�=�>�? P <   �4�4�4�4�4�4�4�4�4555%5/595C5M5O6t6�6l7�<�>�>�>   ` \   x00�0�0�0�0�0�0�0�0 1�1�1�1�23�344�4h5�5�67�7+8�89�9&:�:+;�;K<�<w=�=o>�>[?�?   p 0   ?0�0B1�1[2�2�2�2l7q7�7�7h8m8_;�;g<�<[=�= � H   `2�2�2b7�7�788?8�8�8�8�8�9�9�9O:t:�:�:;x;�;<�<o=�=b>�>w?�?   � 4   o0�0�1�1o2�2H3�3n4H678t8�8�9�9f:�:=;�;<   �    0p89   � p   +2�2K3�3{45�5&6.6�6�6�6�6777R7X7e7�7�7�7�78,8084888<8@8�8�8�899 9<9:H:p:u:�;�;0<5<R=b=�=�=*>�>   � L   �0�0�0�0�0X2p23�3
4o4�4?5�5w6�6�7
888%8�8�8�9�9�9�:;};k>�>K?�?   � L   /0�0+1�1$2�23t3�3[4�4;5�526�6+7n7�7_8�8W9�9R:�:O;�;R<�<b=�=�>?o?�? � 4   M0�01�1�1p2�2P3�3@4�4/5�5�6;7�78�89z9:/; 0    �5\6�6�6 @    �9�<�<�< P     �344p4H5�5�5�5H6�68�= `    k6�6�6�6�6�7 p    f4k4�4�4�89*=�=�>   � `   b0�0�0�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333X3|3�3�3[4�4w5�5g6�6[7�7R8�8R9�<�<.>�?   � �   70;0A0E0K0O0U0Y0_0c0i0m0s0w0}0�0�0�0�0�0�0�0�0�01X1]1g1�1�1�1�1�1�1/2_2�2�2�2�2�3�3�3474L4�4�45%5�5�56�6�6�6�6#7Y7�7�7�7�7�7l8�8�8�8�8�8�8:9S9�9�9�9:b:~:`;�;a>�>�>'?.?~?�?�?�?�?�?�?�? � �   0L0�0�01A1�1�1�12)2�2�2�2>3�3�3�3 4l4w4�4�40555�5�5�5�5�5�5�5666&6+666V6_6h6u6�6�6\7c7�7�78<8p8u8 9#9*9I9O9U9y99�9�9�9�9�9�9:&:8:=:O:�:�:�:�:�;�;�;�;�;�<�<�<�=�=�=">,>u>�><?A?x?}?�?�? � x   �0�0�0�1�1�1�2�2�2)4:4R4c4�7�7 8-82878\8h8�8�8�8�9
:7:<:A:s::�:�:�:�:;1;6;;;<<!<&<=??;?@?E?w?�?�?�?�?�?   � P   0/04090�8�8�89"9'9L9X9�9�9�9�:�:;;;H;T;�;�;�;�=>$>Q>V>[>�>�>�>�>�> � (  D2K2U2y2�2�2�2�2�2�233 3'3_3f3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444"4(4.444:4?4D4J4O4U4^4e4l4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45/565=5`56666%6/686?6E6x6}6�6�6�6�6�67U7�7�783898@8Z8�8999�9;:F:�:�:�;�;�;�;�;�;�;�;�;�;�; <7<G<c<�=�=�=3>;>D>T>`>v>�>�>�>�>�>�>�>�>??9?T?�?�?�?   � �   0_0j0s0{0�0�0�0�0�0�0�0�0�0�01121Q1F3X4]4o4o5x5�5�5�5�5�5�5�5�5�5�56)6F6K6�6�677$7E7e7�7�7�78C8Q8�8�8�8�8�89999+949:9C9H9N9V9\9�9�9�9�9@:J:V:r:�:�:�:�:�:�:�:�:�:�=�=�=�=�=>#>(>??/?�?�?�?�?�?�?   � �   00*0J0v0�0�0�0�0�001<1R1d1�1�1�1�12n2t2�2�2�2�23\3h3�3�3�3�3�3�3�344434D4w4�5�5656A6n6s6x6�6�6�6�6�6�6�6�677i7u7W8c8�8�8�899�9�9�98:=:O:c:�:�:�:�:�:;;0;5;R;W;�;�;�;�;A<p<�<�<=F=}=�=�=!>x>|>�>�>�?�?�?�?  	 �   00D0I0N0[0t0�0�0�0�0H1M1_1�1�1�1�1�1�1�13383=3O3)4G5S5v5�5�5�5�5�5�566.6k6777[7f7C8O8|8�8�8�8�8�8�8�89!9N9S9X9�9;;/;[;`;�;�;<*<U<w<�<�<�<=A=�=�=�=�>�?   	 �   000N0I1l1|1�1�124292>2m2�2�2�2�4�4�4�4�4/5;5h5m5r5%6y7�7�7�78 8M8R8W8�8�8�8�8�8�9<<@<]<�<�<�<=�=�=�=�=�=�>�>�>�>�>�> ????3?    	 �   '0]0l0u0�0�0�0�0�0�0�0111!1+1/191H1L1R1Y1�1�1�1 222)202C2J2�2�2�2�2�233#3(363N3�394?4M4W4�466D6I6N6e6w6�6�6�6�6�6;7G7t7y7~7�7�7�7�7�7�78^8h8�8�8�8x9�9�9�9�9�9�9�:�:�:3;z;�;�;N<U<�=�=�=�=�=�=J>^>�>�>�>�>&?J?Y?n?s?x?�?�?�?   0	 �   a0o0z0�0�0�0�0�0�01U1]1�1!6�6�6�6�6�6T7[7n7�7�7�7�7�7�788878?8H8]8�8^9f9~9�9�98;C;P;X;g;|;�;�;�;�;�;=%=+=?$?l?r?x?~?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @	 �   000$060;0A0G0_0f0�012171<1y1�1�1�1�1-3=3B3H3i344<4C4O4�4�4�4�45]5�5�5A6~6�6�6!7m7�7�7%8q8�8	99e9p9�9�9:(:y:�:�:�:1;};�;�;%<q<�< =x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=`>d>h>l>p>t>x>|>�>�>�>�> P	 8   n1s1x1�1�1�1J2I3N3W4�45�5�6/7�;1<====�?�?�? `	 L   0%000S0^0�044�8�8�8�8(9-9?9W9l9�98:h:�:�:�;�;e<�<
==(=8=D=�>P?�? p	 �   l01;1�1�1�1G2S2�293H3�3�3�34444)4]4m4r4w4|4�4�4�4�4)5.53585B5_5d5i5w5�5�5�6�637�7�7�7�7l8�8�8)9:W:t:�:�:�:�:�:�:;U;#<*<�<�<�=�=�=�=�=�=�=�>�>�>	??1???X?n?�?�?   �	 �   '0-0<0E0N0W0a0u01e1122/2k2t2�2�2�2�2�233333�3�3�344l4u4�4�4�4�4�45�6�6�6�6�6�6F7K7P7X7�7�788'8;8G8b8r8~8�8�8�8�8�8	99%9�9�9�9�9�9�9�9�9 :':�;�;�;�;�;<<<?<H<r<w<|<�<1=J=S=�=�=�=�=�=:>C>L>t>   �	 �    0@0P0U0Z0_0�0�0�0�0K1W1v1�1�1�1�1�1�1�122*2V2r2~2�2�2�2�2)3.333f3k3p3u3�3m5|5�5�5�5�56#606=6U6}6�6�6�6�6�6�67D7[7�7�7�7�8�8�8�8�8�8Q9Z9�9�9�9�9�9::I:N:S:�:�:;1;:;d;i;n;�;�;h=m==�=�=(?-???�?�? �	 $  P0V0\0k0s0{0�0�0�0�0�0�011'161?1Q1n1{1�1�12292L2S2Y2n2t2�2�2�23�3�3�3�344;4L4T4Z4g4�4�4�4�4545>5^5�5�5!6.6<6H6P6�6�7�7�78Y8c8z8�8�8�8�8�8�8�8�89"9(9<9A9I9R9X9l9r9{9�9�9�9:,:d:�:�:�:�:�:�;�;�;<<<<�<�<�<�<�<�<Z=e=�=�=�=�=�=�=�=�=�=	>>(>3>O>Z>�>�>�>�>�>Z?e?t?�?�?�?�?�?   �	   0V1_1|1�1�1�1�1�1�1�1=2L2U2�2�2�2�2�2�2�2�233-3�3�3�3�3�3�3�3�3L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4v7~7�7�7�7�7�7�7�7�7888 8)8=8E8�8�8�8�8$9e9w9�9�9�9�9�9�9�9�9:$:,:x:�:�:�:�:�: ;	;�;�;@<D<H<L<P<y=�=�=�=$>3>9>B>G>k>}>�>�>�>�>�>�><?N?o?|?�?�?�?�?�?�? �	 �   y1�1�1�1�1�1�1�1�12252=2E2M2U2�2�2�2�2�23353=3F3`3n3w3�3*464>4G4P4X4�455*5U5k5s5�5�5�5�5�5�5�5�5�5�56^6}6�6�6�6�6
779788!8*8N8U8o8|8�8�8�8�9:,:Q:a:>;�;�; <<<<<<<< <x<|<�<�<�< �	 $   %1V1o5�57�7�7�7:7;�;�<�=�> �	 x   �0S12�2H3t309I9Q9W9h9z9�9�9�:�;�;�;�;�;�;?<M<U<[<d<j<�<�<�<�<�<�<�<�<�<�<�<==S=[=j=s=y=�=�=�=+?4?>?P?b?m?u?�? �	 �   �1�12282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2�2�2�2�2�283<3@3D3H3L3P3T3X366%6.6M6�67#787d7r7{7�7�7I8Z8i8r8�8�8�9�9�9�9�9�9�9�9:$:-:�:�:�:�:�:;;;�;�;<!<Q<Z<a<�<�<�<�<�<�<===3=<=\=e=l=�=�=�=�=>>1>9>>>�>�>�>�>�>�>�>�>�>�>�> ???  
 @  Y0r0{0�0�0�0�0�0�01'171@1c1k1(2:2e2u2�2�2�2�2�2�2�23�3�3�3�3�3(4�4�4�4�4�4�4�455'595K5X5z5�5�5�5�5�5�5�5�56!636E6X6a6�6�6�6�6�6 77k7r7{7�7�7�7�7~8�8�8�89 9$9(9,9094989<9@9D9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9 ::(:,:�;�;�;<<$<-<2<G<V<e<t<�<�<======= =1>B>a>f>u>�>�>�>�>�>�>�>�>4?8?<?@?D?H?L?P?T?X?�?�? 
 �    00.0<0D0P0\0k0t0�01p1}1�1�1�25*585E5�6�6�6)727@7I7|7�7�7�7�7�7�7�7�788i8w8�8�8�8�8�9�9�9�9~;�;�;�;�;<<<�<
=b=�=�=�=�=`>�>    
 �   I2`2n2w2�2�2�2�2�23;3�3Y4�4z5�697y7g8�8�8�89X9i9�9�9�9�9�9�9
:(:I:W:`:;;�;�;�;�;<�<�<=6=V=v=�=�=�=�=>6>V>v>�>�>�>�>t?   0
    �3�9�9I; @
    ^2�4�5d6�7?<�>? P
 d   60N1v182K2�3F5�5�586D6U6`6i6w6�6�6�6�6�6&7�9X:�:�:�:�:�:9;W;d;�;�;<===�=�=�=�=>>�>�>�? `
 4   �0�0�0�0�0'23�3�4�5�6w7g8W9G:';(?�?�?�?�?�? p
 x   00)020?0�0�0�0C1�1�1�1�122+2Y2�2�2�2�2�2�2�2�2�2$34'4S4c4m4�4�4�4i5�56d6�6757|8�9�9�9�9�9�9�9�:�:<;U;�?�? �
 p   0(0D0`0|0�0�0�01�1�1�1�1�12E2y2�23g4�4O5[5�687=7O7r7�798�9;�<�<�<�<�<==?=D=I=�=�=�=�=�=�=�=>">'> �
 �   70C0	1171<1A1�1�122!2�2�2�283=3B3�5�5�5�5�5�5�5�56?6]6d6h6l6p6t6x6|6�6�6�6�6�6�6B7M7h7o7t7x7|7�7�7�7 88888888f8l8p8t8x8�9�9�9�9�9 ::F:�<====L=U=�=�=�=�=>L>U>>�>�>�>�>�>�>?�?�?   �
 �   E0L0x0�0�02191�1�1�1�1�122F2K2P266s6|6�8�8
9<9T9[9c9h9l9p9�9�9�9�9�9�9�9�9�9�9 :J:P:T:X:\:�:�:�:�:�:�:�:;G;y;�;�;�;�;�;�;�;�;�;�;�;�;�;H>M>_>x>�?�?�?�?�?�? �
 �   �0�0�0�0�0I1R1[1c1�1�1�122"2-292l2s2y2�2�2�2�2�2�2�2�2�2�2�2�2�233i3u3}3�3�34@4G4q4}4�4�4�4�4�4�4�4�45566/6\6h6{6�687=7O7�7�7�7�7�7�7m8y8�8�8�8�8H9[9a9::::: :";5;�;�;�;
<<+<4<^<c<h<�<�<�<�<�<�<==$=V=_={=�=�=�=�=�=�=�=�= �
 `   �2�2�3�3;5G5�5�5,7�7�7�7�7�7f8x8�8�899N9S9X9�9�9�9�9�9�:�:�:Y;e;�;�;�;I<P<^=e=�>�>w?   �
 h   B0�0O1[1�1�1�1p2�2�2"3)3X3_3�8�8�8�8�8�8�8 9999999094989<9@9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9 �
 �   1�1�2�2�2�2�2 3333�3�3�3�3�34 4%4y4�4�4�4�4�4�4555'5.53585B5I5N5S5]5j5o5u5}5�5�5�5�5�5�5�5�5�56*616K6V6]6u6|6q7z7�7�7�7�7�7:8C8m8r8w8�8�8!9J9S9}9�9�9::5:^:g:�:�:�:�:�:j<s<�<�<�<�<�<R=Y=�=�=�=�=�=F>O>�>?2?[?d?�?�?�?�?�?   �
 �   �1�1�1�1�1#2+2j2s2�2�2�2-343a3�3�3�3�3�344Z5c5�5�5�5�5�5<6D6�6�6�6�6�6-767�7�7878@8j8o8t8�8�8�:;);L;"<.<�<�<�<�<�<�>�>Y?a?�?�?�?�?�?�?     �   ?2G2?3G3S4Z4�4�4*525�5�5�5�5:6F6s6x6}6�6�6�6�6�6�8�8(9-929q9z9�9�9�9�9�9�9�:�:�:�:�:�:�:;;;(;7;�;�;�;�;�;�;�<�<�<�<�<�<==)=.=4=A=F=L=�=�=�=>>>>J>V>b>g>l>�>�>�>�>�>�>�>�>#?(?-?2?�?�?�?�?    �   0000=0B0G0�0�0�0�0�0�0�01"1T1�1_2�2�2�2�2�233!3?3D3I3�3�3�5�56�6�6�677/757P7]7b7h7u7z7�7�7�7�72878<8A8t8�8�8�8�8�8�8�89999$9M9R9W9\9�9�9�9�9-:2:7:<:g:l:q:�:�:�:�:;;;.;7;i;�;t<�<�<�<�<�<3=:=I=i=n=s=�=�=*>1>;>M>W>w>|>�>�>�>     �   y1�1�1�1�1�1�1�1�12222"2)2.232=2J2O2U2]2g2n2s2y2�2�2�2�2�2�2
33+363=3U3\3H4Q4{4�4�4�4�45
5535<5f5k5p5�6�6�6�6�6�672777<7�=�?�?   0 0   �0�0�04�4�455(56^6$78/888�8�8�8�8   @ �   �2�2>3q3�3�3�3�3�3�3�3 44X4]4o4�4�4�4�4�455/5o5}5�5�6!7i7�7�9�9�9�9�:;;/;y;�;�;�;�;�;�<�<�<�<>">(>3>9>E>l>?�?�?�? P \   *0/040\3%4�4�4�4q6�6X7�7�7�7�9\:h:�:�:�:�:;";Y;o;�;�;4<J<|=>>>>]?i?n?s?�?�?�?   ` T   	111�1�1�12[2`2e2�2�2�2333�344;4j4�5%6M6�6+7U7�7>�>�>2?�?�?�?�?�?   � 4   �78c8�9�9�9�9�9:!:6:B:n:W<u<�<�<�<W==�=   � D   01�1�1�1�1%2�4�4�4�4535R5q5�5�5�5�56�6�6�6�67,7f7�7�?�?   � X   �0a1m1�1�1�162a3h3�4�4�5�5�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;H;L;P;I>S>w>Y?   � @   Y5�5!7&7+707�7�7�7�7�7�7�7�78!8&8+8_?h?�?�?�?�?�?�?�?   � �    0�1�1�1�1�1p2�2�23_3h3�3�3�3�3�3444�5�5b6n6�6�6�6�6�67 7%7N7�7�7�7�788"8`8g8�9�9�9�9�92:>:k:p:u:�:�:�:k;�;�;2<><k<p<u<�<�<;>�>�>�>�>R?u?~?�?�?�?�?�? � �   0<0A0F0�0�0�0�1262E2x2�2�2�23Q3t3}3�3�3�3�3�3484=4B4{4�4�4�5�5�52676<6b6�6�6�6�6�67F7�7�7�7808G8S8y8�8+9J9�9:#:H:�:�:�:;O;t;�<�<�<�=�=>2?G?�?�?�?   � �   0070�0�3�3�3�3�3�4�451565;5]5�5�5�5�5�5�5�5�56
66"60666f6o6�6�6�6�6]7n7�7�7�7�778X8a8}8�8�8)929\9a9f9�9�9�9�9�9::":)<4<F<]<�<�<�<=/=4=9=�=�=>>>�>�>??5?:??? � �   �1�12!2&2�234�466�6�6�6�6�6(707�7�7�7�7�7]8d8�8 9=9I9v9{9�9!;*;T;Y;^;�;�;�;�;<<#<�<�<�<�<�<$=)=.=�=�=�=�=>2>7><>|>�>   �   K0T0~0�0�0�0�0�0�0�0#1+1n1w1�1�1�1�1�12"2'2�2�2*3/343q5}5�5�5�5�5�5666U6]6�6�6�6�6�6"7.7[7`7e7[8g8�8�8�8):f:o:�:�:�:�;Y<�<�<�>    �   d1p1�1�1�1�1�1V2b2�2�2�2�23�3�3�3�3�3445�5�5�5�5�5686=6B6K8�899K9P9U9�9�9�9�9�9�98:?:�:�:�:�:�:;;I<U<�<�<�<�<�<= =%=g=�=�=!>�>�>�>�>'?,?1?q?y?   �   1m1;2D2n2s2x2�2�2�2�2�233b3k3�3�3�3�3�3444�4�4'5,515�7�7�7�7�7�7�7"8'8,8g8o8�8�8�8�8�869B9o9t9y9x:�:�:�:�:\<�<�<	===U=a=�=�=�=A>v>�>1?8? 0 t   G0N0�1�1f2/3�3b4n4�4�4�4�56666=6k6r6�;�;�; <<<<<<<< <$<(<@<D<H<L<P<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<   @ `   3+3X3]3b3�3�3�3�3�3�5�5(6-626�6707b7�7�7�7�7;8D8n8s8x8�8�89	997>M>�>�>(?9?}?�?�?�?�? P     0&0P0U0Z0�5�5�9�9�=�=z> ` (   222�4�4�4�8�8�8�;�;�;�<�<=   p <   �4�4�4�5�5�5(6-6?6�6�6�6h8x8�8C9	;�;�;�;�;�;r<�>�>   � h   0'030b0p0~0>2L2�2�2>3L3�3�3�6888 8$8�:�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � <    000000�3b405J5�5�5�5�5�5688�8�8D9�:!>'>|>�> � T   �0�0�0.1*2w2�2�2�2�2s3�3�5�5)6�:�;�;<<<�<�<�<=J=V=�=�=�=�=�=>>>b?�?   � �   �0�0�0�0�0�1�1�1�1�142�2�2333�3�3�4	595>5C546@6p6u6z6�7�78"8'89$9T9Y9^9":):�;�;7<C<s<x<}<G=S=�=�=�=�>�>�>�>�>�?�?�?�?�? � �   �0�0111�1�1222�2�3�3444�4�4555�5	6�6�6777�7�788!8�8�8�8�89�9�9*:/:4:�:�:-;2;7;�;�<�<�<�<�<="=�=�=�=�=%>,>�?�?�?�?�?   � x   �0�0�0�0�0�1�1222�2�2$3)3.34'4W4\4a4+575g5l5q5D6P6�6�6�6T7`7�7�7�7{8�8�8�8�8�9�9�9�9�9�:�:�:�:�:�;�;�;�;�;   � t   J1V1�1�1�1>2z3�3�3�3�3 4$4(4,4044484<4@4D4H4L4P4T4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4$5(5,5054585<5@5   � \   6�6�6�6�6�6V7h7�7�788>8C8H8�8�8�8�8�8t9�9�9:2:7:<:�:�:;4;9;>;�;�;�<=8>?>?�?     p   G0�0�0*1/1412�2�2�2�2�2�2�8�8�8�8�8094989<9@9D9H9L9P9T9X9\9`9d9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9  �   H1M1_1�1�1�1E2�2�2�2�2%3+343I3�3�4�4�455"585�5�5�56(646@6V6�67&7^7c7h7�7�7�7�7�7�78�8�8�899�9�9�9�9:K:i:H;M;_;�;�;<<�<�<�<�<�<x=�=�=�=M>V>!?�?   �   �0�0�011.1D1m1z1�1�182=2O2x4}4�4�4�4�4535O5y5�5�5�6�677-777V7�7C8O8�8�8�80999c9h9m9R:�:�:�:;@;l;�;�;<<#<e<q<�<�<�<Q=�=�=�=>>>d>�>�>   0 |   00A1H1%2�2q3!4-4]4b4g4C5�5�5�5�5*616�;�;<	<<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$= @ P   �6�7�7�7�7�78)8Y8^8c8�9�9;;>;C;H;�;�;&<+<0<~<T=[=m>y>�>�>�>�?�?�?�?�? P |   S1_1�1�1�1�2�2�2�2�2�3�355�5�5�5�5�5�6�6�6�6�6A8M8}8�8�8S9_9�9�9�9:@;L;|;�;�;R<^<�<�<�<=�=x>�>�>�>�>�?�?�?�?�?   ` �   k0w0�0�0�0�1�1�1�1�1�2�2�2�2�2�3K4W4�4�4�4�4�4]5d5�5�5�5�5[7g7�7�7�7m8y8�8�8�8�9�9�9�9�9�:�:�:�:�:�;�;<<<�<�<%=*=/=>>>>C>H>? ?P?U?Z?   p �   ;0G0w0|0�0M1Y1�1�1�1c2o2�2�2�2u3�3�3�3�399B9G9L9�9;;N;S;X;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�< � (   (<-<?<e<n<�<�<�<i=�=�=4>@>??   � �    2^2�23^3�3N4�4�5
6.6j6�6�6:7�7�78 8J8O8T8�8�8�8�8�8�:�:�:�:�:�:;';Q;V;[;<<D<I<N<�<�<�<�<�<�< =*=/=4=�>�>�>???D?P?}?�?�?�?�?�?�?�?   � �   �0�0�0�0�0�0�0111L1U11�1�1r2{2�2�2�2�3�3�3�3	44<4A4F4l4�4�4�4�4�4�45!5Z5c5�6�6�6�6�677;7@7E7�;�;==�=�=�?�?�?�? � �   00R0W0\0�0�0�0�0�0�01Q1Z1P2g2�2�2�2<3E3�7�7�7�7�7�7�7�7�788888 8&8,82888>8D8J8P8V8\8b8h8n8t8z8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89
9999"9(9.949:9@9F9L9R9X9^9d9j9p9v9|9�9�9�9�9�9�9�9�9;	; ;Z;�;�;�;< �    O<Y<�<   �    =   � X   1114 4$4(4,4<7@7H8H=L=P=T=X=\=`=d=h=l=p=�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �   111111 1$1(1,1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1,2024282<2@2D2H2L2P2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2445 5$5(5,54585�5�5�5�5�5�5�5�566 6074787<7@7D7H7L7P7T7X7\7`7d7h7l7�:�:�:�:�:�:8?<?@?D?H?       <8@8D8H8L8   0 8   0242,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�? @    �7�7�7H>L>P> P �   H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<   ` ,   �0�0�0�0�0�0�0 111111 1$14181<1 � ,   @0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0   �    t=�=�=�= � �   `4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7 �     x8|8�8�8�8�8�8�8�8�8�8�8 � L  $4(4<4D4H4P4h4t4�4�4�4�4�4�4�4�4�4�455,5D5L5P5X5p5�5�5�5�5�5�5�5�5�5�5�5 660646H6P6X6p6�6�6�6�6�6�6�6�6�6�67777,7D7H7\7`7t7|7�7�7�7�7�7�7�7�788$8,80888P8\8t8�8�8�8�8�8�8�8�8�8 9990989@9X9p9t9�9�9�9�9�9�9�9�9�9�9::0:H:P:d:h:|:�:�:�:�:�:�:�:�:�:�:�:;;4;8;L;T;X;\;d;|;�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>> � $  014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�3�3�3�3444484X4x4�4�4�4�45(545X5x5�5�5�5�5686X6x6�6�6�6�6�6787X7x7�7�7�7�788 8X8t8x8�8�8�8�8�8�89$909h9t9�9�9�9�9�9:$:H:T:`:�:�:�:�:�:;;4;<;H;L;X;l;x;�;�;�;�;�;�;�;<<,<0<L<P<l<p<�<�<�<�<�<�<�<===P=\=�=�=�=�= > >,>P>p>�>�>�>  D   00<0\0|0�0�0�01d1�1�1�1�12@2�2�2�2�2�2�2�2�2�2�243<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444�4�48:@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=H>X>h>x>�>�>�>�>�>�>�>�>�>     H   �0�0�041@1D1H1L1P1T1X1\1`1d1p1t1x1|1�1�1�1�1�1�1�1�1�1�45�8�8�8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    