MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ,gfhs5hs5hs5�H�5is5s��5ss5s��5s5a~�5ks5hr59s5p�5ss5s��5[s5s��5is5s��5is5Richhs5        PE  L z��O        � !
  �  �     �4                             �                              � X     (                            0 4?  `�                                            �! �                          .textbss�                        �  �.text   �     �                   `.rdata  X  �    �             @  @.data   �D   �     �	             @  �.idata  	         �	             @  �.reloc  8J   0  L   �	             @  B                                                                                                                                                                                                                                                                                                                ������F� �/ �I �W� ��( ��� ��e ��� �^g �9� 鴨 �O� �* �%\ �C 髊  �V� �1� � �gX �w � �B �� �  ��W �$� �� �Z0 �@ � h 雺  �& ��u �* �W> �V ��� ��t �j �> ��` �$� �Ye �z� �� �p�  �+ ��  �W �� 駖 颹 ��� �H �7 �9 �	 �m �� �
t �ui �P�  雧 �� ��K ��� �g� ��
 �c �h� ��0 �^. �1 �ą �?�  �:> �E� �� �[R �F� ��� �,T �� �4 �]� �H�  �c� �� 驪  �" ��� �ړ �� �p� �+5 � ��� ��Z ��c �" �m� ���  � �� ��  �Ԋ ��1 �*� �� 進 ��� 閤 �3 �L� �'Z ��� �� �x� �3n �.� ��� �Tn �� ��y  �U�  �? ��J ��  �qY �l 駪  �� �� �
 ��� ���  �ɬ  �t< �: 銰  �e �� � �֘ �qK ��# ��� ��& �� �< 郟 � ��~ �< �? � �Ep �p� � �f�  � �\  ���  �� � �C � � �I� �� �  �
k 酅 �Ђ �o ��� �� �� � ��� �; �x� �J � ��Q �d�  ��  �Z\ �� ��3 �k2 ��a �� �, �'� �a �� ��  �S5 �bc �I$ ��H �� ��  ��s  �$b �$ �f ��F �̐ �GZ  ��f ��3 �W �#�  �^�  �Iv  ��3 �O� �� �%/ �  �h �V �!�  ��  �; �"k �-� ��� �� �^�  �y< �4 � 骫 �U� ��7 �k� �a �j 霟 �� ��= �R 鈿 �C) �- �Y� �$� �O�  �� �� �6 �; �V� ��  �|Q �� 鲸 �=� 阷 � ��  �I� ���  �OH ��S �uv �( �9 �v: �!/ ��� �� 邷 �͟  �� 飬 �a ��k �T � �u �) � & �� ��� �Q ��H �k �b ��[ � �� 龈  �I� ��> �� �*H �U	 �p �+� �6S ��q ��Y  �E �C �m�  �H
 �3� �> �	 �� �o� �� � ���  � �f �� �< �G� �R� �� ��, ��� �>� �h �4O �� ��A �Ũ ��_ ��j �J �� �<�  ��_ �G �}O �X� ��a �Y �y�  �d�  �_i ��  �� �Z �[�  �F` ��� �| ��9 �B� �? �(p  �Ӹ �G �i� 鴳 �5 ��O �5X �P5 �M �&� �qI �8_ �7� �y �]� �� �D �>�  �_ �2 ��� �� ��p ��  �� �6. �Ah �Lu � �bT �; �(� �c �Ε �� �9 �2 �z �" �`i �� �&; �c_ �l�  駑 �b. �} �XM ���  �.�  �	� �% �^ �
� �� ��� �% ���  �1E �,  �e] �RW �m� 騑 �s� �~ �� �4� �o) �� �u � �a^ �� �� �,& �w�  �% �R ��Y  �#� � �v �Dz �O ��< �3 ��V �� ��0 �a< �l% ���  �" �}�  �Ț �#p �n �9�  �T< �? 麪 �v �� 雴 醴 �� �l� �W �� �> �س ��  ��Y �: �� �\ �� ��9 ��� �c ��� �1� �" ��  ��� �� 騂 �D ��� �^b � ��  �o  �\ ��@ �ۋ  �f� � ��� �W2 ��. �]V �H�  �C; �^& �U] �� �� �Z2 �u� � ��4 �� �o  �B �C �r� �m�  �7 ��� �W ��� �D� �?� ��  �yb �p� ��� �6� ��  �K �� �"� �mz �� ��C �r �5 �Ԧ �O" � � �p�  �` ��@ �au �,� 闆 �2� �]� �X� � ��M �	� �T �_� 銸 �U? � ; ���  �" �E �� �� �RD �< �� �C! �~� �T �} �O' ���  � � $ �� 鶡 �� �D �C �B�  �
 �XU �CH ��� �W �vZ �� ��� ��� � �� 醞  �A. �ܔ ��0 ��Y �-� � �Z �  �9 �t� �O� �
� �� �0 �4 �9 �/ ��w �'� �"h �mf �H| �C �� ��{ ��0 �oC �* �T � � � �v �!w �̵  鷣  �� ��� �x� �. �: �� �� �f �� �K � �K� �z �m 鬗  �� �2� �=� ��  ��  �>C �= �d# �� �
 � �Y �k� �f �� �� �Y �� �E � �#� �N; �U �4 �� ��� �3 � � ��: �H �� �d � �� �=c � �S �� �i� �DC �� 銍 �%�  �@w  ��, �fF �# � �7� 颉 �� �XL �S� ��  �  ���  �_o  �*� ��  �p �[ �f 鱦 鬨  ��� �� �=w �V ��% ��  �	�  �D ��' ��, ��" � 1 �e �O �1�  �A �� ��b  �M; �ȟ  �� �nA �i� �d� �9 �J�  �Q � ? 黅 ���  �q� ��� �gm �X �0 鸻 � �� �[ � ��m �d �W �� �r �] ��  �" ��1 �R �-� �� �c' �+ ��� �3 �W �D �? �� �kG �j ���  � �w� �� �m ��  �s�  �>� ��; �. �_� 麺 ��[ �� �+g �6� �� �<G ���  �W � �a �	 �� �� ��V �o ��o �u3 �� ��� �6� �a� �|� �7 ��� ��� �< �< �� �i� �D� �B �+ 酬 �p� � �v �7W ��  �ge �r� �� � �Y ��� �� �$�  �� �k �uw �, �K( �V�  �H �f �KU �B� �� ��� �� �>� ��L ��  �/= �� �u� �`- 鋄 �xV ��� ��< �� �R�  �  ��� �C� �4 ��m �Ľ �O�  �Z�  �� ��O �k �v� ��� �<k ��� �w �mz �h�  鳭 ��X �	 ��{ �� �
_ �U� � � ��� �F�  � �|  闟 �"
 �]� �� �C` �� ��? ��f �< �J
 ��  �  �- 鶄 �r �� �ww ��A �͵ ��  �SN �.k �Y� �4H ��J 隲 �5� �  ��% �V�  �A� �,x �': �? ��� �� �3� �� �� 餈 �' �m �5\ �0� ��� �fs  �M �l� �1= ��� �� �S �SF �.h �� �� ��4 �z� �eq �F �6 ��T �! �,� ��\ �Rx �͖ ��X �S� ��. 陲 鴚 ��� ��  ��� ��  �K�  �6 �� �, �x  �r� 靗 �8� �CH �b �� �4  �?� ��  ��B � � � ��� ��w ��h �w�  �� � �; �S� �I �)� 鴟  �Ol �:� �� �� 黼 �F> �1
 鬦 �	 �� 鍫  �� �3� ��� �y� 锴 �� �� �� ��^ � �� �a� �,� �7�  �"* �m� ��| �T �� �8 ��$ ��c 隶 �, � �f �f4 ��L �� �	 �K �-6 �h�  �- �^� �9 �D�  �u  ��) � �8 ���  �F �R � ���  �B� �- �H� �#� �T �y�  鄂 �� �z� �%Q �`z  鋐 �` ��# 鼱 �7� �� �x �8 飝 �n�  �I �$� �� �z� ��Z � � �kC �F� �1y �3 �Q �� �ݮ �7 �F �3 �? �  �Q �. �E ��u ��  �& �Q �L �7� ��5 ��D �h� 铿 龻 �9�  �3 �/� ��}  �Ź �  �+& �vH �A ��& �7 �Ra �� ��+ ��  �� ���  �t� �Od  ��`  �e� � r  �P 馰 � ��H  �� 鲦 �h �� ��a �P �9� �T% �/� �� �� �� ��I �f} �! �\8 �ǥ �"> �= ��� �� �~� ��1 �	 �� �Jn � �@[  ���  �fC �� �X �P �2� ��D �X� �F �s �0 �D. � ��j �� � � �� �/ �y �, �	 ��� �-z  �H� �W �� ��y �4� 鏀 ��I ��6 �	 �k] �@O �� �O � ��4 �M~ �y �8 �G �	� �n  � �z� �U= �` �|  �f �q� �| �W� �R1 ��$ �� �s�  �ޥ �Y�  �<O �/ �
� �5� �I �[� �f� �Q_ ��� ��T �� �� �� �� �>Y �R ��  ��N �J 鵅 ���  �@ �6� �
 �L� �ע ���  �: �hA �� �Nu  �	 �5 �. �T ��$ �p$ �[� ��; �! �
 �'� �r �  ��� �$ �$ ��# �� �	 ��� �
 ��# �� �&X ��i 鼁 ��$ �B  �=� ��V ��. ��& �Y' ��� �/�  ��� �%� ��\ �;^ �z ��7 �L �'� ��  ���  �X�  � �. �g �D� �� �Z] 鵚 ��" �k� �&� �A� ��" ���  ��% �-� �R ��N  ��{ ��b �$- �O� �3 �e� �P� ��  ��( �A# �" �L �� �mt �h0 ��G �>� �i~ ���  �?Q �� �5\ �0� ��3 �f�  �q�  鬾  �� �b= �� �H� �=M ��V �Y8 ��� �� �� �% ��V �� �&� �� �<N �71 �^  ��: �HL �#�  �^5 �	r �� �/ �5 �� �� �c �f� �A ��| 鷻 �� �� �X� �S� ��n � �M  �K � �5� � �K� �B �A�  �\( �  �"v  �~ �H� �v �� 陴 �x ��� ���  �E�  �p� �۟ 閘 �A�  ��* �2 � �M�  �� �3 �^� ��B 鴭 鏧 �7 �� ��� ��� �F �1?  ��5 ��� �� �]E �� �C� ��
 �9* �=" �� �Z� �� � F  � �ֳ �!� �<w �'< �R� �-� �ȉ �y �^A �	� �� �_[ �jB �E- � � �[	 �� �w �< �'� 鲄 ��V �8� 部 ���  � �t�  �� �Z\ �!I � $ �+� �v� �� ��� 鷤 ��� �=� �(� �c � � �t ��L � 镻 � �  ��� ��t �UJ �,L � ��  ��I �X �#8 ��  �I�  �$� �� � �" ��; ��0 �V� �! �|� �w� �r( �7 �x� �3z ��G � �4� �� �zu � �` �3 �6 �A�  �s 釋 �Rh ��_  �= �� �, �I� �$�  �# � �e  � �  �� 鶠 ��� ��/ �� �� ��|  ��x ��� ��N � �8 �[H �_ ��B  �` ��$ ��  �q�  �* �W: ��x �} ��� �#> �� ��5 �t* �?  �:� ��  � x �K �< �H �L� �g� ��0 �-� �� ��n  �n> �i�  ��q  �G �z� ��� ��p � �� ��� ��D �'u  �b
 ��� ��G �Ӎ �^V �� �, �� �` �u1 ��^ �k �� �ab ���  �wF 钺 �-\ �x} ��, �] � �$G �/� �:� �5< �@+ �[n �F- �aQ �,! �; 颁 �=� ��P ��| �^  �L  �t� ��O �J! �5� �M �� �v5 ��] �� �� ��� �( �� � �N* �� �, ��� �
$ �%5 �` �� �V� �4 �� �7�  ��2 青 �� �c� ��= � �S �_ � �
 �
 ��	 �6� �� � �� �� �M
 ��	 �s  ��  �	�  ��( �� �J^ �$ �0� ��� �
 �� ���  �G �Rh �B �hN �C� �n� �I! ��q �5 �z �% ��$ �{ �V� ��� ��� �7�  钔  �=G �8 鳊 �.� �] �d�  ��D �j� ��� �`6 �{�  �c ��P �� ��B � �}k �[ �3. �~6 �	; �� �@  ��D �%� �0 雓  ��  �A� �m  �W� �R� �m �rD �S, ��1 �	5 �DJ �n �� �%� ��� �5 �R �Q� �\� ��  �� � �� 鳚 ��� � �t �+ �Z �� �; �+� �D �Q �� ��G �"� �M� ��
 �Å ���  �D �xD �?e  �Z� �e ��: �[" �V� ��h �<�  �W� � 靕 �h� 郆 �n� ��  �t� �� �J ��Z �zD ��  ��?  �a+ �,� 鷟  �  �=�  鈏 �� ��. �GC ��Y �/- 麊  �b  �h �;� �& ��� �� �wk �"� �m � �$ �>� ��) �( 鯣 �ʤ  �u' �0� ��3 �! ��  �� � 钇 ��f  �h� �P �~7 �. �r ��  �P �� �PW ��H  ��X �Q) �,�  �g�  �<C �-� �- �C�  ��� �� �B �_n �Z �� ��c �� �� �� �* ��� �u �* �� ��N �w � �TN �- �r �U@ ��� �W ��� � �<�  �R �l ��8 �8� �3 龱 �I �d$ �OC ���  �e% �s �� ��v � �9  �Ǡ �2� �� � �C�  鞬 �Yk �$% 韋 �z�  ��  �� �A �v�  ��$ �|' 鷔 �B� �]� �6 �A �� ���  �DA  ��J �� ��9 � ��@ �k ��S �L� �� �Be �mF  �(;  �)@ �g  �) 鄔 �_F �Z� �� �I �� �f�  �Q� 霭  �G� �U �� �2@ �3 �n� �J �c �o� ��S �U � �+� ��� �Q� �L� ��g ��� �= �� � 鮩 �YR �b �Z 麱  �@ �@D �{� �K �C �� �5� �r� �=�  �b? �� �� ��� �+ �ߺ �
 �U�  �` �� � �1 �8? �! �: ��� �x� �3) �( 鹁 �t �� �j� �%�  � �  �[�  � �A ��� 釩 ��B ��0 �8� 飱 �. �y_ �B �: ��  �h �T � �v� ��� �l{ �� ��� �-� �Ȯ  �C� � �)� �� �� �z �U6 ��  �˼ �F� ��f ���  �GK �L � �C �3% �~ 鉕 �T� �V �Z� � �� �K �v�  ��l  �ܴ � �# �-| ��$ �� �� �yh �C �߅ �� �e�  �0�  �> �v_ ��� �� �G� �� �ݣ �j ��� �no � �Y �_a �>  鵒 �= �| �ֳ ��> �<� 駲 �b� �}O �6 ��� �> �Y! �t �O3 � �j � " 髱 �x �� �H  �� 鲴 �U> �x ��� �^� �i� �>  韯 �� 鵪 �u �Y �� �, �� ��  �R� ��� �� �S� ���  ��  ��� �?� �Z|  �� � " �� �6 �Af �L� �7� ��X �� �� �3S �� �Y� �T� �OD �� �uf  �' ���  �F� �+ �<� �wC 颌 ��� �(0  �Sq �" �y� �TR �
 �:� �� �P�  �� ��2 �Qp  ��< �8 �j 静 �� 鳈 ��� �C �ԉ �� �:< ��k ��; �; �� �Q �<� �g� 鲎 �-| 鸘 �� �N �� ���  �o
 �m ��� � � �k� � �! �} �0 �"� �! �x� �3� �>� �YG �D% ��� �� � �@� �[V �P 鱗 ��:  �� �b ��x �� �� ��H �g  鴥 �5 �� 饞 �g � �� �a� ��m ��" �® �U: �X^ �n  ��.  �y/ �4f  �Od  �
! � �p� �� �& �a�  �l� �w8 ���  ��  �� ��  �@ �Y �� �?� �� �%h �� �ۜ �6�  � 霆  �� �� �]` ��  �� �n� �	� ��  �� �* �: �P� �k� � �a� ��� �G� � ��5 ��� �B ��{ �% �$� �� �
s �� �P�  �v 関 �A! �,Y �9 �bB 靝 ��� �3Z �.|  �y�  �D{  ��  �B �� �Pc  �[Z  ��� ��O  �\D ���  �� �-) ��A �, �� �u ��= � �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E���Ex��M�U;������EE�E��_^[���   ;�������]� �����������������������U����   SVW��@����0   ������=�� t��EP�����;��9���_^[���   ;��)�����]��������������������������������U���   SVW��������   ������j h������������P�g������E������������}� u��  j h��������{���P�E�P�Ĳ������������������������� t�  j h���� ����=���P�������E썍 ���諨���M������j h����P�������P��8���萧����8���Pj�M��F�����8���������P����^���j h|������������P��h����K�����h���Pj�M�������h����S�������������j�������׹��������Pj�M����������������j h���������Y���P�������ݦ��������Pj�M����������������������諧���}� t1�E�P�������q����M�Q������Rj�M����������������+�E�P�������@���������Qj�M��&����������x����M�苨��R��P�}�׬��XZ_^[��   ;��¾����]�   }����   }sc �����������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��Ž����EPj��MQ�U�R����H�Q�҃�;�螽���E�_^[���   ;�苽����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H$�у�;��+����E�_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H0�у�;�苻���E�_^[���   ;��x�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   ��Ѓ�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;�莺��_^[���   ;��~�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M����   ��;�����_^[���   ;��������]� �������������������������������U����   SVW��@����0   �����������   ������ǀ�   MK衰����u3���   _^[���   ;��v�����]�����������������������������U����   SVW��@����0   ������_^[��]������������U���`  SVW�������X   ������E�������������  #�������  tZ������ tB������t�  �������  �u  ��  ���蝟����u3���  �   ��  �   ��  ��  �E�E��E�    �	�E���E�E��M�;�  �E��H�U�<� u��h@��E��H�U��P�Ѩ������th8��E��H�U��P賨������u1j h ������������������P�G������������L����   h��E��H�U��P�d�������u>�E��H�U���    j h �����������������P������������������8h���E��H�U��P��������u�E��H�U���    �    �  ������   �E�E��} u�s�E��x t�hj h�������������������P�M��	�,���P������R�����P������P�=�����������B����������7����������,���3��3�_^[��`  ;�踶����]���������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   ������EP�M��=����EP�M��[����E�P�M�%����M��*����ER��P�$�轣��XZ_^[���   ;�訵����]Ë�   ,�����   8�s ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��%�����E�P�MQ����B�H�у�;������E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M�����P�M�苳���E�_^[���   ;��w�����]� ���������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B<��;�����_^[���   ;��
�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��BL��;�虳��_^[���   ;�艳����]� �����������������������������U���8  SVW��������   �������&����E��E�E�E�P�M�������M�����������ۅ�����]ă��E��$��`���P�M�萚����褶��������ۅ�����]����E��$��x���P�M��������v���������ۅ�����]��E�]����E��$������P�M��c������B���������ۅ�����]����E��$���E��$�������^���P�M��������E��$������P�M�����������������ۅ����ݝt����E�ܝt���������   �g����l���j hT��� ����ٺ���� ���P�������� ����D���j hz0  �>������E��E�]����E��$���E��$�����襳��P�M��+���j h   jjh   ������P������P�	�����P�{�������h���j艤������h���u1���E��$��0���P�M��
���������������ۅ����ݝt���������Q������E��$�����$��H��������P�M������   R��P������XZ_^[��8  ;��ְ����]�   ������   �time �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVWQ��,����5   ������Y�M��E�� �M���$�n������M����A�$ݝ,����T�����ܽ,����-���_^[���   ;��X�����]� ��������������������������������������������U���<  SVW��������   ������E�E��M������E�j jh�  �������̻��Pj jh�  ������跻��P�������Q���P�M�� ����E��������!����}� t�M�� ���j jh�  ������r���Pj jh�  ��$����]���P�� ��������P�M�覔���Eԍ� ����ǫ���}� t�M�覠��j jh�  ��H�������Pj jh�  ��\�������P��8���蝡��P�M��L����Eȍ�8����m����}� t�M��L���j jh�  ������辺��Pj jh�  ������詺��P��p����C���P�M������E���p��������}� t�M�����j jh�  �������d���Pj jh�  �������O���P����������P�M�蘓���E�������蹪���}� t�M�蘟��j jh�  �������
���Pj jh�  ����������P������菠��P�M��>����E��������_����}� t�M��>���j jh�  ��(���谹��Pj jh�  ��<���蛹��P������5���P�M������E�����������}� t�M�����j jh�  ��`����V���Pj jh�  ��t����A���P��P����۟��P�M�芒���E���P���諩���}� t�M�芞��j jh�  �����������Pj jh�  ����������P������聟��P�M��0����E��������Q����}� t�M��0����   _^[��<  ;�踫����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��BL��;�藪��_^[���   ;�自����]������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E��M�H�E�_^[��]� �����������������������U���H  SVWQ��������   ������Y�M��E�E�M�谗���E������$h�  ������P�M��I�����躣���]Ѝ������I��������$h�  ������P�M�������艣���]������������N����E��M�褗���E��E�P�M������M��2���������ۅ�����]����E��$�M��լ��������ۅ����ݝp��������$h�  �M�����ݝ`���j ��@���誢���E������������t�=  �E��4���j ��4����r���� ��(���j ��4����]���� �������(����������������  ��  �������  t�������  ��  ��  j h����������j�M�茓���E�P� �����ǅ���    �������������ۅ���ܝ`���������   �����$������  P�M�� ���ݝ �����݅ ����$��@���肣�����E��$�����P��@����N���݅p���� ���$������蘩��P�M�����j h   jjh   ������P������P�������P�n������������E�P��������  Q�M��8�����tj hz0  蝱����j�P�������������E��$�����$����������P�M�腗��j�M��5����[j�M��)����E���������Dz�����$�E�P����������E��$�E�P�h�����j�M�������E�P�x�����j ��@���蔠��ǅ(���   ��@����g�����(���R��P�|��g���XZ_^[��H  ;��R�����]� ��   ������   ��@���   ��myarray time �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M����   ��;��ɤ��_^[���   ;�蹤����]� �����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B�Ѓ�;��U���E��P�M�Q����B@�H�у�;��3���_^[���   ;��#�����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B�Ѓ�;�赣���M��#���P�U�R����H@�Q�҃�;�萣��_^[���   ;�耣����]� ������������������������������������U����   SVWQ������:   ������Y�M��M��ۉ����E�P�M�Q����B@�H$�у�;��	����E�P�M�נ���M�蝌���ER��P�������XZ_^[���   ;��Ѣ����]� �   �����   �bc ���������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B,�Ѓ�;��E���_^[���   ;��5�����]����������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bt��;��ס��_^[���   ;��ǡ����]������������������������������U����   SVWQ��4����3   ������Y�M��M��i����E��t�E�P詏�����E�_^[���   ;��T�����]� ������������������������U���  SVWQ�������`   ������Y�M��E�E�M�������E��M�襇��h&F �������В��P������賔��j �E�P������Q�M�-����������������.��������� tuh�f �M�薱���E��}� t#j ������赚��Pj�M��L�������������h&F �������L���P�������/���j �E�P������Q�M����������谝��ǅ����   �M�赩��������R��P�̛����XZ_^[�Ā  ;�������]� �   ԛ����   ��d ����������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�M�Q������   �H`�у�;�����_^[���   ;��ޞ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U���P  SVWQ��������   ������Y�M��M豤��P�M�m�����u3���  �M�����E�M裋���E��E�    �M�袄���M�蚄��j jhq  ������迪��P�M�袑���}� tj �E�P�M���������   j��p���P�E�����j h���������g���������Pj��p����d����������ͅ��jj��p������������$j��p���誄��j �������$���P����������������P��p���Q�U�R�M�ͫ��������������������v�����������t8ǅ���   ��p���舆���M��N����M��x����M��p���������  ��p����Z��������$h�  �M�訖������W�����d���ǅX����  ���X�������X�����X���;�d����  �}� ��  �E�   j j��X���P��,����!���P��������������Q�M��7��������舙���}� tj �E�P�M��W�������  j��@���P芁����P�M�������@����y���jj�M��V���jj(�M�����j j'�M�����j h����\����t�����\���Pj�M��t�����\����݃��hq  �������U���P�������8���������P�M�Q�U�R�M�����������w���������誘����w�����t-ǅ����   �M�荘���M�跄���M�评����������  ǅL����  j j��X����L���P������迧��P������蟎��������Q�M��ը���������&���j������P�D�����P�M�轌���������3���hg j�M�����jj�M��ϐ��j h��������7�����L�����X�����y���R������P�n�����P�����Q�� ���R�@�����Pj�M������� ����l����������a���������V�����L�������L���hq  ��T���迋��P��D���袍����D���P�M�Q�U�R�M�k����������;�����D���������;�����t*ǅh���   �M�������M��!����M�������h����Q�E�    �����ǅt���   ��t���P�MQ������ǅ����   �M�褖���M��΂���M��Ƃ��������R��P�آ����XZ_^[��P  ;��������]� �I    �����   *�����    �����   �p���   �maingroupBc cid linkboxBc frameBc ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E�M��E��E_^[��]��������������������������U����   SVW��(����6   �������EP��,���Q����B�H(�у�;�胖��P�M�˟����,�����~���E_^[���   ;��\�����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P0��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P4��;��q���_^[���   ;��a�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M��B,��;�����_^[���   ;��ܔ����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P8��;��q���_^[���   ;��a�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B��;������_^[���   ;�������]������������������������������U���  SVWQ��L����m   ������Y�M��M�v����E�E�P�M�R����M�m�����L���ۅL����]ă��E��$�M�������L���ۅL����]������$h�  �M��K����]��E�    �	�E����E��E��]�������   �����$�E��  P�M������]��EP�M����  Q�M��מ����|����E��E�������Dz6��|��� t-�����P��|����`��������P�M�3w��j j�M�����d���j 貅����3�R��P�d�耀��XZ_^[�Ĵ  ;��k�����]� �I    l�����   �����`   ��m1 time ����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;�莑��_^[���   ;��~�����]� ����������������������������������U���4  SVWQ�������M   ������Y�M�������P����QH�M��B,��;������   ���}�E_^[��4  ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP����QH�M��B0��;�腐��_^[���   ;��u�����]� �������������������������U���,  SVW�������K   ������h'  �)w����P�M��s����M�豙����uǅ����   �M��bx���������   j h�������������j h�������讘��j ������P������������l���P�����Qh=8j	�U�Rh�� 蠇����������������臛���������w����������w���M���w��������R��P����Y}��XZ_^[��,  ;��D�����]Ë�   ������   ��path �������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�輛�������_^[���   ;�蕎����]����������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVW��0����4   ������h��jUh��j裕������8�����8��� t��8�����x����0����
ǅ0���    ��0���_^[���   ;��������]���������������������������������������U����   SVWQ��4����3   ������Y�M��M��@����E�� L��E�_^[���   ;��O�����]����������������������U����   SVWQ��4����3   ������Y�M��M��#z���E��t�E�P�9{�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��\����E�� ���E�_^[���   ;�������]����������������������U����   SVWQ��4����3   ������Y�M��M��ћ��_^[���   ;��+�����]������������������U����   SVWQ��4����3   ������Y�M��M���x��_^[���   ;��ۋ����]������������������U����   SVWQ��4����3   ������Y�M��M��1����E��t�E�P��y�����E�_^[���   ;��t�����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��t���E�� ��E�_^[���   ;�������]����������������������U����   SVWQ��4����3   ������Y�M��M���}��_^[���   ;�車����]������������������U����   SVWQ��4����3   ������Y�M��M��w���E��t�E�P�x�����E�_^[���   ;��T�����]� ������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|.h��h�   h��hp�������h��h�   ��r�����EP�M�����_^[���   ;�踉����]� ��������������������������������������������U����   SVW��@����0   �������EP�MQ����B��0  �у�;��C���_^[���   ;��3�����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|.h��h�   h��hp�������h��h�   ��q�����E��H�U��_^[���   ;�蘈����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@   �M������EP�M��v���E�_^[���   ;��	�����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M�诓��_^[���   ;�談����]������������������U����   SVWQ��4����3   ������Y�M��E��HQ���E�$�M�����_^[���   ;��K�����]� �������������������������������U����   SVWQ������9   ������Y�M��E��8 tD�E�    �E��H�M��E�    ��E���E�M����M��E��M�;H}��E�P�h~�����E��     �E��@    �E��@    �E��@    �E��@    _^[���   ;��v�����]�������������������������������������������������������������U���  SVWQ�������G   ������Y�M��} �M�������   �;  �E��x uh��h�  �	o����3��  �E��H�U�D
��M���y���U��B��E�U��E�    �E�    �E�    �E��x ta�E�    �E�    �E��H�M���E؃��M܃� �E؉M܋Ũ��ŰE��@��������������M�;�����|�U�;�����s븋E��@��������������M�;�����u�U�;�������  �E��M;H~3�E��@��������������M�;������~  �U�;������m  j j�E�P�M�Q��o���E��U��E���������������E�;�����uE�M�;�����u:�E�;E�|2�M�;M�r(�E��������������E�;�����K|�M�;�����s>�   ��t.h��h�  h��hp��I�����h��h�  �Em����3��U  �E��8 u@��h��h�  j j�E�P�M�Q�o��P����B���  �у�;��ԃ���U���D��h��h�  j j�E�P�M�Q��n��P�U��P����Q��  �Ѓ�;�莃���M���E��8 u3��   �E��H�U���ȋU��J�E�M��A�E��HQ�U��R�E��HQ��u�����E�    �E�    �E��H�M���E؃��M܃� �E؉M܋Ũ��ŰE��������������E�;�����#|�M�;�����s�E�Pj�[�����������맋E��M�H�   _^[��  ;�谂����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��} }3��.jjj�EP�M��O�����u3���E��H�U�E�Ѹ   _^[���   ;�������]� �������������������������������U���P  SVWQ�������T   ������Y�M��} }3��  �} 
�   �  �E��H;M~�U��B�������	�M������������U�U�E��x uh��h@  �i����3��3  �E��H��9M��  �E��H+M�U��J�E��x ��  �E��@�؃��M���y���U��B��E܉U��E��@�E�U�j jRP�,k���ẺUЋE̙�������������E�;�����ud�M�;�����uY�E��@�E�U��������������M�;�����|5�U�;�����r(�E��������������E�;�����K|�M�;�����s>�   ��t.h��hO  h��hp��o�����h��hO  �kh����3��  �E��@�E�U��M��A�E��@�E�U��M��A�E��8 u8��h��hV  �E��H��Q����B���  �у�;���~���U���<��h��hW  �E��H��Q�U��P����Q��  �Ѓ�;��~���M���E��8 u3��W  �E��H�U���ȋU��J�} ��   �E��H+M��Q�E��ȋ�+M�u��E���j jVQ�li���U�BP�EE�M��Q��P�v�����E��P�E�+E�U�j jRP�1i���M�AP�U��BP�Rv�����;�E��H��Q�E�+E�U�j jRP��h���U�BP�E��H�U��P�v�����?�} ~%�E��P�M��QR�E��H�U����Q��u�����E��H�U���ȋU��J�  �E��H�U�D
��M���y���U��B��E��U��E��@��������������M�;������~  �U�;������m  j j�E�P�M�Q�/h���E��U��E���������������E�;�����uE�M�;�����u:�E�;E�|2�M�;M�r(�E��������������E�;�����K|�M�;�����s>�   ��t.h��hw  h��hp��}����h��hw  �e����3��*  �E��8 u@��h��h{  j j�E�P�M�Q�fg��P����B���  �у�;��|���U���D��h��h|  j j�E�P�M�Q�&g��P�U��P����Q��  �Ѓ�;���{���M���E��8 u3��  �E��H�U���ȋU��J�E��M��A�E��M;H}2�E��H+M��Q�U��B�M��R�EE�M��Q��P��s�����E�    �E�    �} ti�E��H;M}5�E��H�U��B��Q�U��E+B��P�M��Q�E��H��R�m�����E��H�U��P�M��Q�U��B�M��R�m�����} ��   �E��H;M}M�E��H�M��U��B�M��Q�E���E����E��M����M��E�;E}�E�Pj���������������E�    �E��H�U�щE���E����E��M����M��E�;E}�E�Pj�Ή�����������ЋE��M�H�   _^[��P  ;��#z����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E;Et��EPj �MQ�e����_^[���   ;��x����]�����������������������������������U����   SVWQ��4����3   ������Y�M���j j�����P�M��B��;��w���E�_^[���   ;��w����]��������������������������U����   SVWQ��4����3   ������Y�M���j �EP����Q�M��B��;��Cw���E�_^[���   ;��0w����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EPj�����Q�M��B��;���v���E�_^[���   ;��v����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M��ƃ��_^[���   ;��Kv����]������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;���u��_^[���   ;���u����]���������������������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M�Ck���E�_^[���   ;��u����]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M����   ��;��u��_^[���   ;��u����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;��t��_^[���   ;��t����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;��!t�������_^[���   ;��
t����]� ������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��~����E�M�� f��_^[���   ;��s����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BX�Ѓ�;��2s��_^[���   ;��"s����]�������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;���r��_^[���   ;��r����]� �������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M���Z��_^[���   ;��Nr����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bl��;���q��_^[���   ;���q����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M���Y��_^[���   ;��^q����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��΁���E�EP�M�����_^[���   ;���p����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��p��_^[���   ;��rp����]� ����������������������U����   SVWQ��(����6   ������Y�M���EP����Q�M����   ��;��p���E�}� u3���M��6s��_^[���   ;���o����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B�Ѓ�;��o��_^[���   ;��ro����]�������������������������U����   SVW��<����1   ������} t�E��<��������iU����<�����<���Q�UR�EP��f����_^[���   ;���n����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��X`��_^[���   ;���m����]������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q����B<�H�у�;��mm���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����d��������
ǅ���    �E��@    _^[���   ;���l����]���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��\���E��t�E�P�Z�����E�_^[���   ;��dl����]� ������������������������U����   SVWQ������?   ������Y�M������P�X����P�M��\�������������[�������_^[���   ;���k����]���������������������������U����   SVWQ��$����7   ������Y�M��E��x ufh���t���Ph��j�s������,�����,��� t�MQ��,����u����$����
ǅ$���    �U���$����B�E��x u3��Q�E��x t�E�3Ƀ8 �����9��EP����Q<��Ѓ�;���j���M���E��@   �E�3Ƀ8 ����_^[���   ;���j����]� �����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@   ����H<��Q��;��Cj���M���E�3Ƀ8 ����_^[���   ;��!j����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �4�E��x u3��'��E��HQ�U��P����Q<�B�Ѓ�;��i��_^[���   ;��i����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u����H��#��EP�M��R����H<�Q�҃�;���h��_^[���   ;���h����]� ��������������������������������U����   SVW��@����0   ���������[��_^[���   ;��h����]���������������������U����   SVW��@����0   ������EP����Sx��_^[���   ;��:h����]�����������������U���  SVW�������B   ������EP����x��P�M��Bq��j hL�������p��j �E�P�����Q�M���l�������������������P����������t�M�Im���M���O���E�9j�E�P�M��g\��j�j��EP�M�Q�M��qf���E�P�M�p���M��O���ER��P����MU��XZ_^[��  ;��8g����]Ë�   ������   ������   ��str pos ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��uf���E�_^[���   ;��bf����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��B@��;���e��_^[���   ;���e����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PH��;��e��_^[���   ;��qe����]� �������������������������������������U���,  SVW�������K   ������EP����#u��P�M��bn��j hL���������m��j �E�P������Q�M��j��������������������0M����������t�M�ij���M��M���E�   j�E�P�M��Y��j�j��EP�M�Q�M��c��j hL�������Tm��j �E�P�����Q�M��i�������������������L����������t�M��i���M��L���E�9j�E�P�M��Y��j�j��EP�M�Q�M��c���E�P�M�Qm���M��VL���ER��P�����Q��XZ_^[��,  ;���c����]Ë�    �����   �����   �str pos ����������������������������������������������������������������������������������������������������������������U���P  SVW�������T   ������EP����s��P�M��Rl��j hL���������k��j �E�P������Q�M���g�������������������� K����������t�M�Yh���M��K���E�>  j�E�P�M��tW��j�j��EP�M�Q�M��~a��j hL��������Dk��j �E�P������Q�M��yg��������������������J����������t�M��g���M��J���E�   j�E�P�M���V��j�j��EP�M�Q�M���`��j hL��������j��j �E�P�����Q�M���f�������������������J����������t�M�Qg���M���I���E�9j�E�P�M��oV��j�j��EP�M�Q�M��y`���E�P�M�j���M���I���ER��P����UO��XZ_^[��P  ;��@a����]Ë�   ������   ������   ��str pos ��������������������������������������������������������������������������������������������������������������������������������������������U���t  SVW�������]   ������EP����cp��P�M��i��j hL��������i��j �E�P������Q�M��Me��������������������pH����������t�M�e���M��UH���E��  j�E�P�M���T��j�j��EP�M�Q�M���^��j hL��������h��j �E�P������Q�M���d���������������������G����������t�M�%e���M���G���E�>  j�E�P�M��@T��j�j��EP�M�Q�M��J^��j hL��������h��j �E�P������Q�M��Ed��������������������hG����������t�M�d���M��MG���E�   j�E�P�M��S��j�j��EP�M�Q�M���]��j hL�������g��j �E�P�����Q�M���c��������������������F����������t�M�d���M���F���E�9j�E�P�M��;S��j�j��EP�M�Q�M��E]���E�P�M�g���M��F���ER��P����!L��XZ_^[��t  ;��^����]Ë�   ������   ������   ��str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������EP����Q<�B�Ѓ�;���\��_^[���   ;���\����]���������������������������������U���p  SVW�������\   ������ǅ����    j h���������Ue��P�H�����E���������D���}� u3���   �E�    �E�P�M��|M���E�P�M�Q�M��\������   �}���   �M��L���E��}� tF�EP�������a��������Pj������Q�M���b������������F����tǅ����   �
ǅ����    ��������������������t���������������C����������t���������������C����������t�EԉE�������E�R��P����UI��XZ_^[��p  ;��@[����]Ë�   ������   ������   ������   ��browse dat id ��������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��=B�������_^[���   ;��@Z����]� ��������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;���Y��_^[���   ;���Y����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BT�Ѓ�;��rY��_^[���   ;��bY����]�������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R����P�M����   ��;���X��P�M�@b���� ����BA���E_^[���   ;���X����]� �������������������������������������U���d  SVW�������Y   ������ǅ����    �} u6j h���������?a��P��C�����E�������@���} u3��$  �E�    �EP�M��fI���E�P�M�Q�M��oX������   �}���   �M��~H���Eă}� tF�EP�������]��������Pj������Q�M���^������������B����tǅ����   �
ǅ����    ��������������������t���������������?����������t���������������?����������t�E��E��2�+�}�u%�}� t�EP�M��}@�����.B����t�E��E��������E�R��P����E��XZ_^[��d  ;���V����]ÍI    ������   �����   �����   ��browse dat id ��������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BH�Ѓ�;���U��_^[���   ;���U����]�������������������������U����   SVW������:   ������} u3��   �EP�M���F���E�    �E�    �E�P�M�Q�M���U����tT�}�t�}�u"�EP�M���E��P�{G������t�   �*�$�}�u�EP�M��q>�����"@����t�   ��3�R��P����C��XZ_^[���   ;���T����]�   ������   �����   �����    �dat id browse ����������������������������������������������������������������������������������U����   SVW��@����0   ���������H<��Q��;��2T��_^[���   ;��"T����]�������������������������U����   SVW��@����0   ������E������� _^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��5Y����E�P����Q$�BD�Ѓ�;��mS���E�_^[���   ;��ZS����]���������������������������������U����   SVWQ��4����3   ������Y�M��M��X����E�P����Q$�BD�Ѓ�;���R����EP�M�Q����B$�Hd�у�;���R���E�_^[���   ;��R����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��X����E�P����Q$�BD�Ѓ�;��=R����EP�M�Q����B$�H�у�;��R���E�_^[���   ;��R����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��UW����E�P����Q$�BD�Ѓ�;��Q����E�P�MQ����B$�HL�у�;��kQ���E�_^[���   ;��XQ����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�BH�Ѓ�;���P���M��;9��_^[���   ;���P����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HL�у�;��aP��_^[���   ;��QP����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q$�M��B��;���O��_^[���   ;���O����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP����Q$�M��Bl��;��eO��_^[���   ;��UO����]� �������������������������U����   SVWQ��4����3   ������Y�M�����P$��M��Bp��;���N��_^[���   ;���N����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B�Ѓ�;��N��_^[���   ;��uN����]����������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q����B$�H�у�;��N��P�M�VW���� ����X6���E_^[���   ;���M����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H�у�;��qM��_^[���   ;��aM����]� �������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H �у�;���L��P�M�V��������m<���E_^[���   ;���L����]� �������������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H$�у�;��NL��P�M�V���������;���E_^[���   ;��'L����]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M���A������3��������A;���E_^[���   ;��K����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B(�Ѓ�;��5K��_^[���   ;��%K����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�Bh�Ѓ�;���J��_^[���   ;��J����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H,�у�;��QJ��_^[���   ;��AJ����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H0�у�;���I��_^[���   ;���I����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H4�у�;��QI��_^[���   ;��AI����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H8�у�;���H��_^[���   ;���H����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B$�HL�у�;��QH���E�_^[���   ;��>H����]� ����������������������������������U����   SVW������9   ������EP�M��Q����EP�M�Q����B$�H@�у�;���G���E�P�M�}Q���M��I7���ER��P�8��5��XZ_^[���   ;��G����]�   @�����   L�fn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H@�у�;��G���E�_^[���   ;���F����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H<�у�;��F��_^[���   ;��qF����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H<�у�;��F�������_^[���   ;���E����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H$�QP�҃�;��~E��_^[���   ;��nE����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HT�у�;��E��_^[���   ;���D����]� �������������������������������������U����   SVW��@����0   ���������H$��QX��;��D��_^[���   ;��D����]�������������������������U����   SVW��@����0   �������EP����Q$�B\�Ѓ�;��*D��_^[���   ;��D����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q$�B`�Ѓ�;��C��_^[���   ;��C����]� �����������������������������U����   SVW��@����0   ���������H(����;��CC��_^[���   ;��3C����]��������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;���B���E�     _^[���   ;��B����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR����P(�M��B��;��BB��_^[���   ;��2B����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B��;���A��_^[���   ;��A����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B��;��UA��_^[���   ;��EA����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B��;���@��_^[���   ;���@����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P ��;��a@��_^[���   ;��Q@����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ����B(�M��P��;���?��_^[���   ;���?����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B$��;��^?��_^[���   ;��N?����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B(��;���>��_^[���   ;���>����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B,��;��z>��_^[���   ;��j>����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B0��;��
>��_^[���   ;���=����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B4��;��=��_^[���   ;��=����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BX��;��%=��_^[���   ;��=����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B\��;��<��_^[���   ;��<����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B`��;��E<��_^[���   ;��5<����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bd��;���;��_^[���   ;���;����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bh��;��e;��_^[���   ;��U;����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bx��;���:��_^[���   ;���:����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bl��;��:��_^[���   ;��u:����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bt��;��:��_^[���   ;��:����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bp��;��9��_^[���   ;��9����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��,����t2�M��Q�M��x,����t�U��R�M��e,����tǅ0���   �
ǅ0���    ��0���_^[���   ;���8����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��C����t8�MQ�A�$�M��qC����t"�UQ�B�$�M��[C����tǅ0���   �
ǅ0���    ��0���_^[���   ;��68����]� ������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��77����t2�M��Q�M��$7����t�U��R�M��7����tǅ0���   �
ǅ0���    ��0���_^[���   ;��7����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M��(����t<�M���A�$�M���'����t$�U���B�$�M���'����tǅ0���   �
ǅ0���    ��0���_^[���   ;���6����]� ����������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��1����tE�M��Q�M���0����t2�U��R�M���0����t�E��$P�M���0����tǅ0���   �
ǅ0���    ��0���_^[���   ;���5����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��C.����tE�M��Q�M��0.����t2�U��R�M��.����t�E��$P�M��
.����tǅ0���   �
ǅ0���    ��0���_^[���   ;��5����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��m����tE�M��Q�M��Z����t2�U��0R�M��G����t�E��HP�M��4����tǅ0���   �
ǅ0���    ��0���_^[���   ;��N4����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��|?����tE�M��Q�M��i?����t2�U��0R�M��V?����t�E��HP�M��C?����tǅ0���   �
ǅ0���    ��0���_^[���   ;��~3����]� ��������������������������������������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M�������u3���   �}� u)������8��P�M���������7���   �   ��hP��x���P�M�Q����B���   �у�;��2���E��}� uj��M��3��3��Lj �E�P�M�Q�M������u�E�P�*����3��&j �E��P�M�Q�M�34���E�P��)�����   R��P��	�1 ��XZ_^[���   ;��2����]�    �	����   �	����   �	c len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B�H�у�;��Q1���E�_^[���   ;��>1����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;���0��_^[���   ;��0����]� �����������������������������U����   SVWQ������?   ������Y�M��M��6���E�P�M���(����uǅ���    �M����������$�E�P�M���ǅ���   �M���������R��P�����XZ_^[���   ;���/����]�    �����   �str ��������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�P�M��N!����u3���E�����؋M��   R��P���O��XZ_^[���   ;��:/����]� ��   �����   �c ��������������������������������������U����   SVWQ��4����3   ������Y�M��} ����Q�M��9��_^[���   ;��.����]� ��������������������U����   SVWQ������=   ������Y�M�j �M�%�����E���hP��|���P�M�Q����B���   �у�;��4.���Eԃ}� uj��M��4/��3��dj �E�P�M�Q�M�2���E�P�M�������t �M�Q�U�R�M���5����tǅ���   �
ǅ���    ������E�E�P�m%�����E�R��P�4���XZ_^[���   ;��-����]�    <����   Hmem ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;���,��_^[���   ;���,����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bh��;��n,��_^[���   ;��^,����]� ����������������������������������U����   SVWQ������<   ������Y�M��� ���P�M�!��P�M��08��������� ����H�������_^[���   ;���+����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B8��;��d+��_^[���   ;��T+����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B<��;���*��_^[���   ;���*����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B@��;��*��_^[���   ;��t*����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��BD��;��*��_^[���   ;��*����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BH��;��)��_^[���   ;��)����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P|��;��1)��_^[���   ;��!)����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BL��;��(��_^[���   ;��(����]� �������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P(�M��BT��;��A(��_^[���   ;��1(����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P(�M��BP��;���'��_^[���   ;��'����]� �����������������������U����   SVW��@����0   ���������H(��Q��;��b'��_^[���   ;��R'����]�������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;���&���E�     _^[���   ;���&����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP����Q(�M����   ��;��N&��_^[���   ;��>&����]�( ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B(�H�у�;���%��_^[���   ;��%����]���������������������������������U����   SVW��@����0   ���������H,��Q,��;��b%��_^[���   ;��R%����]�������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B4��;���$��_^[���   ;���$����]���������������������������������U����   SVW��@����0   �������E�Q����B,�H0�у�;��$���E�     _^[���   ;��o$����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B8��;��
$��_^[���   ;���#����]���������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B<��;��#��P�M�H-�����������E_^[���   ;��k#����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q����B,�M��P@��;���"��P�M�F,���� ����H���E_^[���   ;���"����]� �������������������������������������������U����   SVW��@����0   �������j j ����H,��҃�;��l"��_^[���   ;��\"����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H,�Q�҃�;���!��_^[���   ;���!����]� ����������������������������������U����   SVW��@����0   �������E�Q����B,�H�у�;��x!���E�     _^[���   ;��_!����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;��� ��_^[���   ;��� ����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�� ��_^[���   ;��z ����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�� ��_^[���   ;��
 ����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B ��;����_^[���   ;������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B$��;��:��_^[���   ;��*����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B(��;�����_^[���   ;������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B,�M��P��;��Q��_^[���   ;��A����]� �������������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B��;�����P�M�'��������Q���E_^[���   ;������]� �������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��D  �҃�;��@��_^[���   ;��0����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��H  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;��g��_^[���   ;��W����]������������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;����_^[���   ;��s����]��������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;����_^[���   ;������]�����������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;��6��_^[���   ;��&����]�����������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;��Z��_^[���   ;��J����]���������������������������������U���  SVW�������E   ������E�P�M�T���M��������uǅ����    �M��q���������   j�E�P�y������u*�E�P�������uǅ����    �M��2���������Tj�EP�=������u*�EP�������uǅ���    �M�����������ǅ���   �M����������R��P��#�7��XZ_^[��  ;��"����]�   �#����   �#parent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP����Q�B �Ѓ�;��z��_^[���   ;��j����]���������������������������������U����   SVW��@����0   �������EP�MQ����B�H(�у�;����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��  �у�;����_^[���   ;��w����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;�� ��_^[���   ;������]�����������������������U����   SVW������9   ������� ���P����Q�B$�Ѓ�;����P�M�m���� ����6���E_^[���   ;������]���������������������������������������U����   SVW������9   ������� ���P����Q���  �Ѓ�;��$��P�M������ �������E_^[���   ;�������]������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;����_^[���   ;������]��������������������������U���$  SVW�������I   ������ǅ8���    �=� t!������P���{����8��������������������8���������������������������R�M�����8�����t��8����������W����8�����t��8�����������:���E_^[��$  ;������]�����������������������������������������������������������U����   SVW������9   �������EP�� ���Q����B���  �у�;����P�M������ �������E_^[���   ;�������]��������������������������������U����   SVW��@����0   ������j�EP�f�����E_^[���   ;������]������������������������������U����   SVW��@����0   ���������H���   ��;��/��_^[���   ;������]����������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;������E�     _^[���   ;������]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����;��:��_^[���   ;��*����]� ������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;�����_^[���   ;������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��W��_^[���   ;��G����]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B`��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;��u��_^[���   ;��e����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bh��;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bl��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bp��;��%��_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��B��_^[���   ;��2����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��b��_^[���   ;��R����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B|��;���
��_^[���   ;���
����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��
��_^[���   ;��r
����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��
��_^[���   ;��
����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��	��_^[���   ;��	����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��2	��_^[���   ;��"	����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��R��_^[���   ;��B����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��r��_^[���   ;��b����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q����B �H$�у�;��+����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR����H �QL�҃�;��~��_^[���   ;��n����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q����B �H(�у�;������   _^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;��t��_^[���   ;��d����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;����_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;����_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;��$��_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;�� ��_^[���   ;�� ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;��E ��_^[���   ;��5 ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P\��;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B ��;��Q���_^[���   ;��A�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P�M��B$��;������_^[���   ;��������]� �����������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B(��;��a���_^[���   ;��Q�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B,��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B0��;��u���_^[���   ;��e�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B4��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B8��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B<��;��%���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B@��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BD��;��E���_^[���   ;��5�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BH��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BL��;��e���_^[���   ;��U�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BP��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;��v���_^[���   ;��f�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BT��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;�����_^[���   ;��~�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�����_^[���   ;��������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�����_^[���   ;��v�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PX��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��"���_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��B���_^[���   ;��2�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��W���_^[���   ;��G�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��g���_^[���   ;��W�����]������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;�����_^[���   ;��w�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���   �у�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;�����_^[���   ;��{�����]����������������������������������U����   SVW��(����6   �������EP�MQ��,���R����H���  �҃�;�����P�M�U�����,����W����E_^[���   ;��������]���������������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��s���_^[���   ;��c�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�HD�у�;�����_^[���   ;��������]� �������������������������������������U����   SVW��@����0   ���������H8��Q<��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������E�Q����B8�H@�у�;��(����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   ���������H8����;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q����B8�H�у�;��H����E�     _^[���   ;��/�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q�҃�;��>���_^[���   ;��.�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q8�B�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H �у�;��Q���_^[���   ;��A�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q$�҃�;������_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P����Q8�B�Ѓ�;��-���_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q(�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B,�Ѓ�;��)���_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q�҃�;��"���_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q0�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B4�Ѓ�;�����_^[���   ;��	�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H8�у�;�����_^[���   ;�������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��x  �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP�MQ����B��|  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��3���_^[���   ;��#�����]��������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��W���_^[���   ;��G�����]������������������������������U����   SVW��@����0   �������EP����Q�B,�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��(����6   ������M��:�����E�P����Q�B8�Ѓ�;��r����E�P�M�����M������ER��P��W�O���XZ_^[���   ;��:�����]�   �W����   �Wstr ����������������������������������������U����   SVW��@����0   ���������H��Q<��;������_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ����B�H@�у�;��V���_^[���   ;��F�����]�����������������������������U����   SVW��@����0   ���������H��QD��;������_^[���   ;��������]�������������������������U����   SVW��@����0   ���������H��QH��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ�UR����H�QL�҃�;��#���_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B�HP�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP����Q��<  �Ѓ�;��G���_^[���   ;��7�����]������������������������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP����Q���   �Ѓ�;��@���_^[���   ;��0�����]���������������������������������������U����   SVW��@����0   ���������H�􋑼   ��;������_^[���   ;�������]����������������������U����   SVW��@����0   ���������H���  ��;��o���_^[���   ;��_�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�.  ����B���   �у�;������_^[���   ;��������]�����������������������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;��z���_^[���   ;��j�����]���������������������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW������<   ������EPj h��������{���P�M�Q������������������E�P����Q�B�Ѓ�;��l����M������R��P��^�X���XZ_^[���   ;��C�����]Ð   �^����   �^s ��������������������������������������������������U����   SVW��@����0   �������EP����Q�BT�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q�BX�Ѓ�;��J���_^[���   ;��:�����]���������������������������������U����   SVW��@����0   �������EP����Q�B\�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   ���������H��Q`��;��r���_^[���   ;��b�����]�������������������������U����   SVW��@����0   ���������H��Qd��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   ���������H��Qh��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP����Q�Bl�Ѓ�;��J���_^[���   ;��:�����]���������������������������������U����   SVW��@����0   �������EP����Q�Bp�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Qt�҃�;��c���_^[���   ;��S�����]��������������������������U����   SVW��@����0   �������EP����Q��D  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��  �Ѓ�;��{���_^[���   ;��k�����]����������������������������������U����   SVW��@����0   �������EP�MQ����B�Hx�у�;�����_^[���   ;��������]�����������������������������U����   SVW��@����0   �������EP�MQ����B��@  �у�;�����_^[���   ;�������]��������������������������U����   SVW������9   ������M�������E�P�MQ����B�H|�у�;������E�P�M������M������ER��P��d�����XZ_^[���   ;��������]�   �d����   �dfn �����������������������������������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;��S���_^[���   ;��C�����]��������������������������U����   SVW��@����0   �������EP�MQ����B��h  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��d  �Ѓ�;��k���_^[���   ;��[�����]����������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   ���������H�􋑄   ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;��#���_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP����Q��   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;��@���_^[���   ;��0�����]�����������������������U����   SVW��$����7   ������M�蠹����E�P����Q���   �Ѓ�;�������E�P�M�����M��c����ER��P�4i����XZ_^[���   ;�������]Ð   <i����   Hibc �����������������������������������������������������U����   SVW��@����0   ���������H��`  ��;�����_^[���   ;��������]����������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW�� ����8   �������EP��$���Q����B���   �у�;��0����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��������]�����������������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;��s�����]��������������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ����B���   �у�;�����_^[���   ;��������]����������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;�����_^[���   ;��p�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;�����_^[���   ;�� �����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��0���_^[���   ;�� �����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;��P���_^[���   ;��@�����]�����������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;��s���_^[���   ;��c�����]��������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��'���_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;�������u3���E�R��P�Pq菸��XZ_^[���   ;��z�����]�   Xq����   �q����   �q����   |qdata sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;�������u3���E�R��P�@r蟷��XZ_^[���   ;�������]�   Hr����   xr����   qr����   lrdata sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;��������u3���E�R��P�0s诶��XZ_^[���   ;�������]�   8s����   hs����   as����   \sdata sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�	���P�U�R����H0���   �҃�(;��J���_^[���   ;��:�����]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�*���P�U�R����H0���   �҃�(;��Z���_^[���   ;��J�����]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q0���   �Ѓ�(;��n���_^[���   ;��^�����]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;��b���_^[���   ;��R�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H0���   �҃�;������_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;��b���_^[���   ;��R�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;������_^[���   ;��������]�������������������������U����   SVW��@����0   ���������H0�􋑤   ��;�����_^[���   ;��o�����]����������������������U����   SVW��@����0   �������E�Q����B0���   �у�;������E�     _^[���   ;��������]�����������������������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP����Q��T  �Ѓ�;��'���_^[���   ;�������]������������������������������U����   SVW��@����0   ���������H��p  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   ���������H���  ��;��_���_^[���   ;��O�����]����������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�臿��_^[���   ;��w�����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;�蛾��_^[���   ;�苾����]����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���  �у�;�����_^[���   ;�������]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P����Q��X  �Ѓ�;�蘽��P�M�ڽ����,��������E_^[���   ;��q�����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q������   �H�у�;������E�_^[���   ;��ּ����]� ������������������������������������������U����   SVW������=   ������j hLGOg������?���PhicMC�E�P����������������M��ʬ����u�M������M�������E��M�詬��P�M�����M������ER��P������XZ_^[���   ;��������]Ð   �����   �dat ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;��c���_^[���   ;��S�����]��������������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW������9   ������EP��MQ�� ���R����H��t  �҃�;��}�����蓢���� ���������E_^[���   ;��X�����]�������������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;�����P�M�8�����,����:����E_^[���   ;��ɹ����]��������������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;��`���P�M������,���誡���E_^[���   ;��9�����]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��׸��_^[���   ;��Ǹ����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��g���_^[���   ;��W�����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B���  �у� ;��k���_^[���   ;��[�����]����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR����H���  �҃�$;��ض��_^[���   ;��ȶ����]�������������������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q����B��t  �у�;��R���P�M蚿����,���蜞���E_^[���   ;��+�����]����������������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q����B���  �у�;�贵��P�M�������,����-����E_^[���   ;�荵����]������������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;��'���_^[���   ;�������]������������������������������U����  SVW��(����6  ��������3ŉE��E�E�E�P�MQh   ������R�e�����������Ph������Q��4  �Ѓ�;�胴���E�    R��P�|��p���XZ_^[�M�3���������  ;��Q�����]ÍI    ������   ��t ��������������������������������������������������������������U����   SVW��4����3   ������} 3��^�EP�MQ�UR�EP�¯�����E��}� |�E��9E�|/�}� }h�������P诜�����EE�@� �E���E��E�_^[���   ;��`�����]���������������������������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;������P�M�<�����,����>����E_^[���   ;��Ͳ����]������������������������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;��d���P�M謻����,���讚���E_^[���   ;��=�����]������������������������������������U����   SVW������=   ������������u�\h���M�詢���EPh���M��`����EPh���M��O���j �E�PhicMC�����Q������������&����M��9���R��P�\�腟��XZ_^[���   ;��p�����]Ë�   d�����   p�msg ������������������������������������������������������������U����   SVW������=   ������������u�M葶���E�^h!���M�螡���EPh!���M��U���j �E�PhicMC�����Q�������������P�M��������������M��/����ER��P�h��x���XZ_^[���   ;��c�����]Ð   p�����   |�msg ����������������������������������������������������������������U����   SVW������=   �������o�����u�M聵���E�^h����M�莠���EPh����M��E���j �E�PhicMC�����Q���������ט��P�M�۸������������M������ER��P�x��h���XZ_^[���   ;��S�����]Ð   ������   ��msg ����������������������������������������������������������������U���   SVW�� ����@   �������_�����u3��^h#���M�臟���EPh#���M��>���j �E�PhicMC�����Q�ݲ�������B������������������M����������R��P����a���XZ_^[��   ;��L�����]Ë�   ������   ��msg ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B8�Ѓ�;�貭��_^[���   ;�袭����]�������������������������U���   SVW�� ����@   ������������u3��^hs���M������EPhs���M��Ψ��j �E�PhicMC�����Q�m��������Һ������������蘶���M�論�������R��P�������XZ_^[��   ;��ܬ����]Ë�   ������   �msg ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;��4���_^[���   ;��$�����]���������������������������U����   SVW��@����0   �������EP�MQ�UR����H��@  �҃�;������_^[���   ;�谫����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;��D���_^[���   ;��4�����]���������������������������U����   SVW��@����0   ������E�8 t#��E�Q����B��D  �у�;��ͪ���E�     _^[���   ;�贪����]���������������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;��W���_^[���   ;��G�����]������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;�����_^[���   ;��ש����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��P  �҃�;��p���_^[���   ;��`�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��T  �҃�;�� ���_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��X  �҃�;�萨��_^[���   ;�耨����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��\  �҃�;�� ���_^[���   ;�������]�����������������������U����   SVW��@����0   ���������H��d  ��;�迧��_^[���   ;�诧����]����������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q��h  �Ѓ�;��?���_^[���   ;��/�����]��������������������������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;��æ��_^[���   ;�賦����]��������������������������U����   SVW��@����0   ���������H�􋑄  ��;��_���_^[���   ;��O�����]����������������������U����   SVW��$����7   �������EP��(���Q����B���  �у�;�����P�M�������(���脏���E_^[���   ;��ɥ����]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��g���_^[���   ;��W�����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�胤��_^[���   ;��s�����]��������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�蠣��_^[���   ;�萣����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��0���_^[���   ;�� �����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;�谢����]�����������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��W���_^[���   ;��G�����]������������������������������U����   SVW��@����0   �������EP�MQ����B��$  �у�;�����_^[���   ;��ӡ����]��������������������������U����   SVW��@����0   �������EP����Q��(  �Ѓ�;��w���_^[���   ;��g�����]������������������������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   ���������H��0  ��;�蟠��_^[���   ;�菠����]����������������������U����   SVW��@����0   ���������H��<  ��;��?���_^[���   ;��/�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;��˟��_^[���   ;�軟����]����������������������������������U����   SVW��@����0   ���������H���  ��;��_���_^[���   ;��O�����]����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;��������]�����������������������U����   SVW��4����3   ������j �M�����E��}� t�E�P褟�����E�P�.�����R��P�p��q���XZ_^[���   ;��\�����]Ë�   x�����   ��c ������������������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B��  �у� ;�軝��_^[���   ;�諝����]����������������������������������U����   SVW��@����0   ���������H��P  ��;��O���_^[���   ;��?�����]����������������������U����   SVWQ��4����3   ������Y�M��E���P������_^[���   ;�������]���������������������������U����   SVW��@����0   �������EP������   ���   �Ѓ�;�脜��_^[���   ;��t�����]���������������������������U����   SVW��@����0   ���������HL���   ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������E�Q����B@�H�у�;�踛���E�     _^[���   ;�蟛����]��������������������������������������U����   SVW��@����0   ���������HL����;��C���_^[���   ;��3�����]��������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��ؚ���E�     _^[���   ;�迚����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;��R���_^[���   ;��B�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL���   �҃�;��ۙ��_^[���   ;��˙����]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����QL���   �Ѓ�;��b����E�}� u)��j �EP�M�Q����BL���   �у�;��2�����M�蜉��P�M� ���_^[���   ;�������]� ���������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BH��;�蒘��_^[���   ;�肘����]� ����������������������U����   SVWQ��4����3   ������Y�M�������   ��M��BP��;��'���_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��(  �Ѓ�;�貗��_^[���   ;�袗����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��,  �҃�;��;���_^[���   ;��+�����]� �������������������������������U����   SVW��@����0   ���������HL��Q��;��Җ��_^[���   ;������]�������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��h����E�     _^[���   ;��O�����]��������������������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL�Q�҃�;��ە��P�M謓��������o���E_^[���   ;�贕����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��>���_^[���   ;��.�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q�҃�;�辔��_^[���   ;�讔����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��E���_^[���   ;��5�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��Փ��_^[���   ;��œ����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��e���_^[���   ;��U�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B �Ѓ�;�����_^[���   ;��ْ����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��4  �у�;��n���_^[���   ;��^�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B$�Ѓ�;�����_^[���   ;��ّ����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL�H(�у�;��e���_^[���   ;��U�����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B,�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B0�Ѓ�;�腐��_^[���   ;��u�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��  �҃�;�����_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;�蒏��_^[���   ;�肏����]�������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL��  �҃�;�����P�M����������x���E_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B4�Ѓ�;�腎��_^[���   ;��u�����]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P����QL�B8�Ѓ�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�融��_^[���   ;�莍����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�螌��_^[���   ;�莌����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�螋��_^[���   ;�莋����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;�袊��_^[���   ;�蒊����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;��2���_^[���   ;��"�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;����_^[���   ;�貉����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�H<�у�;��Q���_^[���   ;��A�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��Ո��_^[���   ;��ň����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q@�҃�;��^���_^[���   ;��N�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HD�у�;��߇��_^[���   ;��χ����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HH�у�;��_���_^[���   ;��O�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HD�у�;��߆��_^[���   ;��φ����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HH�у�;��_���_^[���   ;��O�����]� �����������������������������������U���,  SVWQ�������K   ������Y�M��M��l��h�  ��������w��P�������y��j �E�P������Q�M��.m��������������������(�����������tǅ���    �M��"����������M��;���������M����������R��P�|��es��XZ_^[��,  ;��P�����]Ë�   ������   ��dat ����������������������������������������������������������������������������U���  SVWQ�������B   ������Y�M�j��������~��h�  ��$����v��P������ox��j������P�����Q�M��Ms����������������������_^[��  ;��\�����]���������������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������}��h�  ��$�����u��P������w��j������Q�����R�M��r��������+����������7���_^[��  ;�蚃����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H(�у�;������E�_^[���   ;��������]� ��������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������{��h�  ��$����jt��P������Mv��j������Q�����R�M��+q������������������׋��_^[��  ;��:�����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M��h��h�  ������s��P�������u��j �E�P������Q�M��i������������������������������t�M������M������E��M��s��P�M� ����M������ER��P����Jo��XZ_^[��  ;��5�����]� �   ������   ��dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BL�Ѓ�;�蒀��_^[���   ;�肀����]�������������������������U���  SVWQ�������E   ������Y�M��M���f��h�  ������r��P��������s��j �E�P������Q�M��ng��������������������h}����������t�M�Z����M��d����E��M��eq��P�M耉���M��F����ER��P�8��m��XZ_^[��  ;������]� �   @�����   L�dat ����������������������������������������������������������������U���4  SVWQ�������M   ������Y�M��M��e��h�  ��������p��P��������r��j �E�P������Q�M��>f��������������������8|����������t��ݝ ����M��4���݅ �����M���z��ݝ����M�����݅���R��P�h��wl��XZ_^[��4  ;��b~����]�   p�����   |�dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B<�Ѓ�;���}��_^[���   ;��}����]�������������������������U���,  SVWQ�������K   ������Y�M��M��d��h�  �������Ao��P�������$q��j �E�P������Q�M��d�������������������z���������tǅ����    �M�蒆����������M�諊��������M��t��������R��P����j��XZ_^[��,  ;���|����]Ë�   �����    �dat ����������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M���b��h�  ������n��P��������o��j �E�P������Q�M��^c��������������������Xy����������t�M脀���M��T����E�,�M��M���M���P�Q�P�Q�@�A�M��&����ER��P�X��i��XZ_^[��  ;��u{����]� �   `�����   l�dat ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�����E����X�E�_^[��]���������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BP�Ѓ�;��z��_^[���   ;��rz����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;��z��_^[���   ;��z����]�������������������������U����   SVWQ������9   ������Y�M���j�EP�M�Q�� ���R����HL���   �҃�;��y���M���P�Q�P�Q�@�A�E_^[���   ;��jy����]� ����������������������������������������������U����   SVWQ������9   ������Y�M���j �EP�M�Q�� ���R����HL���   �҃�;���x���M���P�Q�P�Q�@�A�E_^[���   ;��x����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M��_��h�  ������1j��P�������l��j �E�P������Q�M��_��������������������u����������t�M�|���M�脁���E�,�M��}{���M���P�Q�P�Q�@�A�M��V����ER��P�(��e��XZ_^[��  ;��w����]� �   0�����   <�dat ����������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M���]��h�  �������h��P��������j��j �E�P������Q�M��N^��������������������Ht����������t�M�t{���M��D����E�,�M��=z���M���P�Q�P�Q�@�A�M������ER��P�h��zd��XZ_^[��  ;��ev����]� �   p�����   |�dat ����������������������������������������������������������������U���  SVWQ�������E   ������Y�M��M��\��h�  ������g��P�������i��j �E�P������Q�M��]��������������������s����������t�M�4z���M�����E�,�M���x���M���P�Q�P�Q�@�A�M���~���ER��P����:c��XZ_^[��  ;��%u����]� �   ������   ��dat ����������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M��F[��h�  �������qf��P�������Th��j �E�P������Q�M���[���������������������q����������tǅ���    �M���}���������M��ہ��������M��}�������R��P����b��XZ_^[��,  ;���s����]Ë�   ������   ��dat ����������������������������������������������������������������������������U���  SVWQ�������B   ������Y�M����E�$��������t��h�  ��$����%e��P������g��j������P�����Q�M���a��������p���������|��_^[��  ;���r����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�X�E�_^[��]� �������������������������������U���  SVWQ�������B   ������Y�M��EP�������l��h�  ��$����
d��P�������e��j������Q�����R�M���`��������ko���������w{��_^[��  ;���q����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U���  SVWQ�������B   ������Y�M��EP�������i��h�  ��$�����b��P�������d��j������Q�����R�M��_��������Kn���������Wz��_^[��  ;��p����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H,�у�;��+p���E�_^[���   ;��p����]� ��������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������g��h�  ��$����a��P������mc��j������Q�����R�M��K^���������l����������x��_^[��  ;��Zo����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP��������f��h�  ��$�����`��P������b��j������Q�����R�M��]��������+l���������7x��_^[��  ;��n����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������<f��h�  ��$����
`��P�������a��j������Q�����R�M���\��������kk���������ww��_^[��  ;���m����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������g��h�  ��$����J_��P������-a��j������Q�����R�M��\��������j���������v��_^[��  ;��m����]� ����������������������������������������������U���  SVWQ�������E   ������Y�M��M��fS��h�  ������^��P�������t`��j �E�P������Q�M���S���������������������i����������t�M�q���M���u���E�,�M���o���M���P�Q�P�Q�@�A�M��u���ER��P����Z��XZ_^[��  ;��l����]� �   ������   ��dat ����������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M��&R��h�  �������Q]��P�������4_��j �E�P������Q�M��R��������������������h����������tǅ���    �M��t���������M��x��������M��t�������R��P�����X��XZ_^[��,  ;���j����]Ë�   �����   �dat ����������������������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��M���P��h�  �������\��P��������]��j �E�P������Q�M��nQ��������������������hg����������tǅ���    �M��bs���������M��{w��������M��Ds�������R��P�<��W��XZ_^[��,  ;��i����]Ë�   D�����   P�dat ����������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M���s���E�}�t�}�t�}�tǅ$���    �
ǅ$���   ��$���_^[���   ;��h����]���������������������������������U���  SVWQ�������B   ������Y�M��EP�������l`��h�  ��$����:Z��P������\��j������Q�����R�M���V��������e���������q��_^[��  ;��
h����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������	b��h�  ��$����zY��P������][��j������Q�����R�M��;V���������d����������p��_^[��  ;��Jg����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������Ia��h�  ��$����X��P������Z��j������Q�����R�M��{U��������d���������'p��_^[��  ;��f����]� ����������������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��f��_^[���   ;��f����]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��e��_^[���   ;��e����]������������������������������U����   SVW��@����0   ���������H�􋑘   ��;��?e��_^[���   ;��/e����]����������������������U����   SVW��@����0   ���������H�􋑜   ��;���d��_^[���   ;���d����]����������������������U����   SVW��@����0   �������E�Q����B���   �у�;��ud���E�     _^[���   ;��\d����]�����������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;���c��_^[���   ;���c����]������������������������������U����   SVW��4����3   �������N^���E��}� u3��_��EP�MQ�UR�E�P����Q���  �Ѓ�;��ic����u+�}� t��E�P����Q@�B�Ѓ�;��Ac���E�    �E�_^[���   ;��'c����]����������������������������������������������U����   SVW��@����0   �������EPj �MQ�S^����P�UR�EP����Q���  �Ѓ�;��b��_^[���   ;��b����]���������������������������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���   �Ѓ�;���a��_^[���   ;���a����]����������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q���   �Ѓ�;��Oa��_^[���   ;��?a����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BL�Ѓ�;���`��_^[���   ;���`����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BP�Ѓ�;��e`��_^[���   ;��U`����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�QT�҃�;���_��_^[���   ;���_����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��  �у�;��n_��_^[���   ;��^_����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;���^��_^[���   ;���^����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BX�Ѓ�;��u^��_^[���   ;��e^����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B\�Ѓ�;���]��_^[���   ;���]����]� �����������������������������U���T  SVWQ�������U   ������Y�M��IX���E�}� u3��  �E�    �E�    �E�    �M��!D���M��=H���E�E��E��E��EPh]  �M��S��j j �E�P�M��&F����u��   �M���B���E���E��Eȃ}� ��   �M��"l���E��EȉE��E�Ph�   �sJ������u�   �}� u�~j �M���A���Eԃ}� u�i�E�P�M���L���E�P��_�����}� t��E�P����Q@�B�Ѓ�;��\���E�    �`����E쉅�����M��a���M��F���������W�}� t��E�P����Q@�B�Ѓ�;��A\���E�    �E�P�L_����ǅ����    �M��Xa���M��E��������R��P����J��XZ_^[��T  ;���[����]� �   ������   �����    �cd ctr �����������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;��[Z��_^[���   ;��KZ����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;���Y��_^[���   ;���Y����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B<��;��bY��_^[���   ;��RY����]� ����������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B(��;���X��_^[���   ;���X����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B`�Ѓ�;��X��_^[���   ;��uX����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bd�Ѓ�;��X��_^[���   ;��X����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�Hh�у�;��W��_^[���   ;��W����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��D  �Ѓ�;��"W��_^[���   ;��W����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bl�Ѓ�;��V��_^[���   ;��V����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��>V��_^[���   ;��.V����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M$�H��h��hP�h��h���E��HQ�U R�EP�MQ���E�$�UR�E��HQ�U�R����HL���   �҃�4;��vU��_^[���   ;��fU����]�  ������������������������������������������U����   SVW��@����0   ������E���M���;��U��_^[���   ;���T����]��������������������������U����   SVW��@����0   �������EP�M��M�B��;��T��_^[���   ;��T����]���������������������U����   SVW��@����0   �������EP�MQ�U��M�P��;��:T��_^[���   ;��*T����]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�M��M�B��;���S��_^[���   ;��S����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;��RS��_^[���   ;��BS����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL��   �Ѓ�;���R��_^[���   ;���R����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ����BL�M���H  ��;��RR��_^[���   ;��BR����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M�����PL��M���L  ��;���Q��_^[���   ;���Q����]������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���P  ��;��bQ��_^[���   ;��RQ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���T  ��;���P��_^[���   ;���P����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HL���   �҃�;��oP��_^[���   ;��_P����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL���   �Ѓ�;���O��_^[���   ;���O����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL��   �у�;��bO��_^[���   ;��RO����]� ��������������������������������������U���  SVW�������B   ������M���9���M��aT���} t�M���8����u"ǅ����   �M��,3���M��T���������Qj�M��8��P�M��I���M��8���E�E�E��E�Ph=���<����������M���2���M��S�������R��P�x��g<��XZ_^[��  ;��RN����]�   ������   ������   ��active mu ������������������������������������������������������������������������������U���  SVW�������B   ������M��8���M��S���} t�M��y7����u"ǅ����   �M���1���M��R���������Qj�M��I7��P�M�uH���M��87���E�E�E��E�Ph<���:����������M��1���M��eR�������R��P����;��XZ_^[��  ;��M����]�   ������   ������   ��active mu ������������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����HL���   �҃�;��@L��_^[���   ;��0L����]�����������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;���K��_^[���   ;���K����]��������������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;��cK��_^[���   ;��SK����]��������������������������U����   SVW��@����0   ���������HL��  ��;���J��_^[���   ;���J����]����������������������U����   SVW��@����0   ���������HL��@  ��;��J��_^[���   ;��J����]����������������������U����   SVWQ��(����6   ������Y�M�j\�f   ���E�}� t	�E�x\ u���EP�M�Q�U�B\�Ѓ�;��J��_^[���   ;��	J����]� �����������������������������U����   SVW��@����0   ������h���EPh^� ��Y����_^[���   ;��I����]�������������������������U����   SVWQ��4����3   ������Y�M��7���M���E�_^[���   ;��FI����]�����������������������������U����   SVW��@����0   �����������   �􋑈   ��;���H��_^[���   ;���H����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�P�K�����E��     _^[���   ;��nH����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��(��]����z	�(��]���]����Au	���]�E��������$�7�����E���E����X�M��`E���E�_^[���   ;��xG����]� ��������������������������������������������U����   SVWQ�� ����8   ������Y�M����]����Azǅ$���   �
ǅ$���    ���]����Azǅ ���   �
ǅ ���    ��$���3�;� ������M���E�$��.����������$�6�����E�����E�$�.����������$�]6�����E��X�E����X����Auh8������P�z/�����E����X�}� u�E�� ���M���M��D���E�_^[���   ;��F����]� ��������������������������������������������������������������������������������U����   SVW��@����0   ��������E�$��M����_^[���   ;��E����]������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X�E����X����Auh8������P�>.�����E����X_^[���   ;���D����]� ���������������������������������U����   SVWQ��,����5   ������Y�M����]����Auh8������P�-�������]�E�� �M���$�W4�����M����A�$ݝ,����=4����ܽ,������$�)4�����U�����E�$�4�����E��X�M���A��_^[���   ;��D����]� ��������������������������������������������������������U���0  SVWQ�������L   ������Y�M��E���� �$�+�����]�E����@�$�+�����]�����]�����At����]�����Au�E�����E����X�U  ����]�����Auz����]�����Auj�E���7���E��E���7���E��}� u�E�����E����X�8�E���}��U��E��E��E��E��}� u��E��E��8�M���E��E��x�M��Y��   ���E��$���E��$�C�����=���]����]�����Au.�E��M��]��E��M��]؋E�� �M��M���E��@�M��M��Y���]�����Au���]؋E����X���E��$���E��$�M�����]��E��]��E��]�����]�����A{ǋE�� �u�M���E��@�u�M��Y_^[��0  ;���A����]������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������E�]����Au�E��E_^[��]�����������������������U����   SVWQ��0����4   ������Y�M��E�M��;t3���   �E�x uN�E�8 uF�E�x u=�E��x u�M��9 u�U��z uǅ0���   �
ǅ0���    ��0����   �R�E��x uI�E��8 uA�E��x u8�E�x u�M�9 u�U�z uǅ0���   �
ǅ0���    ��0����M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� �������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��0�������_^[���   ;��@?����]� ��������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M��>���8 t��E�_^[���   ;���>����]����������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M��>���8 t(�E�P�M�>��P�M�Q�M���=�����LK����t�뾃} t�E�M��}� ~�E�P�M���=���8 uǅ$���   �
ǅ$���    ��$���_^[���   ;���=����]� �����������������������������������������������������������U����   SVW��4����3   ������j�k   ���E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;��H=��_^[���   ;��8=����]�������������������������������U����   SVW��@����0   ������h���EPhD � M����_^[���   ;���<����]�������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u���E�P�M�Q\�҃�;��]<���E�_^[���   ;��J<����]���������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;���;���EP�M���I���E�_^[���   ;��;����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��-;���EP�M��:,���E�_^[���   ;��;����]� ����������������������������������U����   SVWQ������;   ������Y�M�j\�������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;��:���EP������d,��P�M��+���E�_^[���   ;��b:����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;���9���EP�M���*���EP�M��Z'���E�_^[���   ;��9����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;��-9���EP�M��:*���EP�M��&���EP�M��&���E�_^[���   ;���8����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�������E�}� t	�E�x` u���E�P�M�Q`�҃�;��m8��_^[���   ;��]8����]������������������������������������U����   SVWQ��(����6   ������Y�M�jd��������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;���7��_^[���   ;���7����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jh�f������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;��I7��_^[���   ;��97����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jl��������E�}� t	�E�xl u���E�P�M�Ql�҃�;��6��_^[���   ;��6����]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��6��_^[���   ;��6����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��~5��_^[���   ;��n5����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u� ����EP�M�Q�U�Bp�Ѓ�;���4��_^[���   ;���4����]� ����������������������������������������U����   SVWQ������:   ������Y�M�jt�f������E�}� t	�E�xt uh ��M�/(���E�:��EP�M�Q�����R�E�Ht�у�;��24��P�M�""��������1���E_^[���   ;��4����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�������E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;��v3���E�_^[���   ;��c3����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jx��������E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;���2��_^[���   ;���2����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�V������E�}� t	�E�x| u�   �#��E�P�MQ�U�B|�Ѓ�;��42�������_^[���   ;��2����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��4����3   ������j�{������E��}� t	�E��x u3���E���H��;��g1��_^[���   ;��W1����]������������������������������U����   SVW��4����3   ������E�8 u�?j��������E��}� t	�E��x u�!��EP�M��Q�҃�;���0���E�     _^[���   ;��0����]��������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j�L������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;��)0��_^[���   ;��0����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��/��_^[���   ;��w/����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;���.��_^[���   ;���.����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �f������E�}� t	�E�x  u3����E�P�M�Q �҃�;��K.��_^[���   ;��;.����]����������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;��-��_^[���   ;��-����]����������������������������������U����   SVWQ��(����6   ������Y�M�j(�F������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;��-��_^[���   ;��-����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;��,��_^[���   ;��s,����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;���+��_^[���   ;���+����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j4�f������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��K+��_^[���   ;��;+����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8��������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;��*��_^[���   ;��*����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�&������E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;��	*��_^[���   ;���)����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jD�������E�}� t	�E�xD u3����E�P�M�QD�҃�;��{)��_^[���   ;��k)����]����������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� u���EP�M�Q�U�BH�Ѓ�;���(��_^[���   ;���(����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jL�v������E�}� u3����EP�M�Q�U�BL�Ѓ�;��`(��_^[���   ;��P(����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�jP��������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;���'��_^[���   ;��'����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�V������E�}� u3����E�P�M�QT�҃�;��D'��_^[���   ;��4'����]���������������������������U����   SVWQ��(����6   ������Y�M�jX��������E�}� u���EP�M�Q�U�BX�Ѓ�;���&��_^[���   ;��&����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;��&��_^[���   ;��
&����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��r%��_^[���   ;��b%����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;���$��_^[���   ;���$����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��J$��_^[���   ;��:$����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��#��_^[���   ;��#����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��$#��_^[���   ;��#����]� ����������������������������������������U����   SVW������9   ������h�   �������E��}� u�M�T(���E�9��EP�� ���Q�U����   �Ѓ�;��"��P�M��+���� �����
���E_^[���   ;��\"����]���������������������������������������������������U����   SVWQ������?   ������Y�M�h�   ��������E�}� t�E샸�    uj ��������P�M����E�9��EP�����Q�U�M����   ��;��!��P�M������������E_^[���   ;��}!����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��� ��_^[���   ;��� ����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3����EP�U�M����   ��;��2 ��_^[���   ;��" ����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;����_^[���   ;������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����E�M����   ��;��V��_^[���   ;��F����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;����_^[���   ;������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u���EP�U�M����   ��;����_^[���   ;�������]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��Z��_^[���   ;��J����]� ����������������������������������������������U����   SVWQ������9   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�M����   ��;�����E��E�_^[���   ;������]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E��     �E��@    �E��@   �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��} u�4�} t�EP�M�O+��� �} t�EP�M�����E�P�M���_^[���   ;������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B@��;��"��_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BD��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bd��;��E��_^[���   ;��5����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bh��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pl��;��a��_^[���   ;��Q����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pp��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;��_��_^[���   ;��O����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bt��;��j��_^[���   ;��Z����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bx��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��B|��;����_^[���   ;��u����]� �������������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bt��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;��2��_^[���   ;��"����]� ����������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;�����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;��R��_^[���   ;��B����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q@�M����   ��;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;��[��_^[���   ;��K����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����Q@�B�Ѓ�;��e���E�E�#Et�E��#E�E��	�E�E�E��E�P�M�Q����B@�H�у�;��"��_^[���   ;������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�HL�у�;��1��_^[���   ;��!����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�BH�Ѓ�;����_^[���   ;������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q@�B�Ѓ�;��9��_^[���   ;��)����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H�у�;�����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H@�Q�҃�;��>��_^[���   ;��.����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H �у�;�����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;��>��_^[���   ;��.����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B ��;��;��_^[���   ;��+����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP������   �M����   ��;����_^[���   ;������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M���D  ��;��(��_^[���   ;������]� ����������������������������U����   SVWQ��4����3   ������Y�M���E P���E�$�MQ�UR�EP�MQ������   �M����   ��;��
��_^[���   ;��
����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ������   �M����   ��;���	��_^[���   ;���	����]� �����������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B$��;��	��_^[���   ;��w	����]������������������������������U����   SVW��@����0   ���������H@��Q0��;��"	��_^[���   ;��	����]�������������������������U����   SVW��@����0   �������j�EPj ����Q@�B4�Ѓ�;����_^[���   ;������]�����������������������������U����   SVW��@����0   �������j�EPh   @����Q@�B4�Ѓ�;��C��_^[���   ;��3����]��������������������������U����   SVW��@����0   �������EP�MQj ����B@�H4�у�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   ���������H|����;��s��_^[���   ;��c����]��������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H�у�;�� ���E�     _^[���   ;�������]������������������������������U����   SVW��@����0   ���������H|��Q ��;����_^[���   ;������]�������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H(�у�;�� ���E�     _^[���   ;������]������������������������������U����   SVW��@����0   ���������H@��Q0��;����_^[���   ;������]�������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;��@���E�     _^[���   ;��'����]������������������������������U����   SVW��@����0   �������EP����Q@���   �Ѓ�;�����_^[���   ;������]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;��P���E�     _^[���   ;��7����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��d  �у�;��^��_^[���   ;��N����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q �BH�Ѓ�;�����_^[���   ;�������]�������������������������������������U����   SVW��4����3   ������}qF t�1�E�E��}� u�#�EP�M��O����E�P�MQ�M�.������B��_^[���   ;��<����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��Pp��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��BT��;��Z��_^[���   ;��J����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��BX��;��� ��_^[���   ;��� ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��P\��;��q ��_^[���   ;��a ����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��B`��;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP�MQ����B��T  �у�;�����_^[���   ;��s�����]��������������������������U����   SVW��@����0   ������h��hE  �M�����������Ph��hE  �M����������P����H��T  �҃�;������_^[���   ;��������]�����������������������������������������������U����   SVW��@����0   ������E�8 t��E�Q����B��у�;��a����E�     _^[���   ;��H�����]�������������������������������U����   SVW��@����0   �������hﾭޡ���H��@  �҃�;������_^[���   ;��������]������������������������������U����   SVW��@����0   ������} t!��EP����Q��@  �Ѓ�;��q���_^[���   ;��a�����]������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   ���������H��   ��;��/���_^[���   ;�������]����������������������U����   SVW��@����0   ������} t�E�x��u�   �3�_^[��]��������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��L����j�EP�I   ��_^[���   ;��,�����]���������������������������������������������������U����   SVW��4����3   ������}s�E   �E��P�������E��}� u3��:�} t�E��Pj �M�Q�������E�� �����E����E���   �E�_^[���   ;��e�����]��������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;�������j�EP�������_^[���   ;�������]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;������j�EP�	�����_^[���   ;��������]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��L����j�EP�I�����_^[���   ;��,�����]���������������������������������������������������U����   SVW��4����3   ������} tF�E�E��=� t�E�x��u�E��P��������E�P����Q��Ѓ�;�����_^[���   ;��|�����]�����������������������������������U����   SVW��4����3   ������} tF�E�E��=� t�E�x��u�E��P���������E�P����Q��Ѓ�;������_^[���   ;��������]�����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��{���_^[���   ;��k�����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;�����_^[���   ;��������]����������������������������������U����   SVW��<����1   ������=�� tI�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;��h����j�EP�e�����_^[���   ;��H�����]�����������������������������������������������U����   SVW��<����1   ������=�� ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;������[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���  �Ѓ�;��S�����EP�MQ�N�����_^[���   ;��1�����]������������������������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� t0��EP�MQ�UR����H���   �҃�;�������0����j�EP��������0�����0����M��E���th�������
P�p������E�_^[���   ;��4�����]�����������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� to�} t0��EP�MQ�UR����H���   �҃�;�������0����.��EP�MQ�UR����H���  �҃�;��d�����0�����0����E��j�EP�R������E��E���th�������P�M������E�_^[���   ;�������]������������������������������������������������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;�����_^[���   ;��{�����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��;���_^[���   ;��+�����]����������������������������������U����   SVW��@����0   �������EP����Qp��Ѓ�;������_^[���   ;�������]����������������������������������U����   SVW��@����0   �������h   ����Hp��҃�;��[���_^[���   ;��K�����]����������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����Bp�H�у�;�������E�     _^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����Hp�Q�҃�;��^���_^[���   ;��N�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����Hp�Q�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����Hp�Q�҃�;��^���_^[���   ;��N�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����Bp�H�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s   ���E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��>���_^[���   ;��.�����]� ����������������������������������U����   SVW��@����0   ������h��EPh�f ������_^[���   ;��������]�������������������������U����   SVWQ������<   ������Y�M�h�   �s������E�}� t�E샸�    u�M�����E�9��EP�����Q�U�M����   ��;��2���P�M�t�������������E_^[���   ;�������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��n���_^[���   ;��^�����]� ����������������������������������U����   SVWQ������<   ������Y�M�h�   �������E�}� t�E샸�    u�M�����E�9��EP�����Q�U�M����   ��;������P�M����������;����E_^[���   ;�������]� �����������������������������������������������U����   SVW������:   ������EP�M������EP�������E܃}� t��E�P�U܋E܋H �RL��;������E�P�M������M������ER��P��R�����XZ_^[���   ;��������]Ë�    S����   Sbc �������������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@�?�E�@8+'�E�@<'�E�@@�K�E�@D�9�E�@H[8�E�@L�7�E�@P�)�E�@l�8�E�@XV8�E�@\_9�E�@`�9�E�@d�8�E�@T�8�E�@h,�E�@pK9�E�@t�8�E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������������U���h  SVW�������Z   ������j h�   ��\���P�[�����j �EP�MQ�UR�EP��\���Q��������E �E�h�   ��\���P�MQ�URj������R��P�0Y����XZ_^[��h  ;�������]Ë�   8Y\����   DYnp ���������������������������������������������������������U����   SVW��@����0   ������EP�M���   Q�UR�������_^[���   ;��������]���������������������U���  SVWQ��\����i   ������Y�M�� ����M���E��8 u��   �EP��l�������j h��������d���P����������j j���l���Q������R������P�������P������Q�������P�����R�������P�E�������������؈�c�������������������������������������������������K�����l����u�����c�����t�E�P��������E�_^[�Ĥ  ;�������]� ��������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP��������M���E�_^[���   ;�������]� �������������������U����   SVWQ��4����3   ������Y�M��E�P�������_^[���   ;�������]�����������������������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����  SVW������z   ������M�G�����tj �EP�MQ��������u3��Sj h   ������P��������EP�M Q�UR�EP������Q�   ��h   ������P�MQ�URj������R��P��^�3���XZ_^[���  ;�������]�   �^����   �^np �������������������������������������������������������������U����   SVW��@����0   ������j �EP�MQ�UR�EP�MQ�z������Eǀ�   #�Eǀ�   �!�Eǀ�   �"_^[���   ;��S�����]�����������������������������������������̋�`L����������̋�`D����������̋�`H�����������U����   SVWQ��4����3   ������Y�M��E�� ��E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��y����E��t�E�P�������E�_^[���   ;��T�����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �_^[��]��������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;�����������
ǅ���    �E�    _^[���   ;��c�����]������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���  ��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���(  ��;�����_^[���   ;��w�����]������������������������������U����   SVWQ������<   ������Y�M������P����Q�M���   ��;�����P�M���������������E_^[���   ;��������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���$  ��;��w���_^[���   ;��g�����]������������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;�����_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   ���������H��  ��;��/���_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ����B��x  �у�;��S���_^[���   ;��C�����]��������������������������U����   SVW��@����0   �������EP����Q��|  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;��r����E�}� u3���EP�MQ�M�����_^[���   ;��E�����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;��R����E�}� u3���EP�MQ�M�����_^[���   ;��%�����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q8�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q����B�H�у�;��%����U��B�E�_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q����B�H�у�;������U��B_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��E��HQ�UR�EP�M��R����H�Q�҃�;������M��A�   _^[���   ;��������]� ���������������������������������U����   SVW��<����1   ������E��<�����<���t��E� ��E���   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$�<l�   �]  �$����$��=$���   �EP�������=�.  }
������&  �} u
������  h ������Ph��j�9������� ����� ��� t�� ��������������
ǅ���    ��������=� t�EP�������   �   �EP�MQ� �������u����   �   �|�����u�$����$�u\�ͼ���|����=� t?����8�����8�����,�����,��� tj��,�������������
ǅ���    ��    �   ����_^[���   ;�������]Ð�j�k�k�j$l�k����������������������������������������������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M���EP����Q�M��Bd��;������E�}� u3��s��hp������P�M��Q����B���   �у�;��v����E��}� u3��4��EP�M��Q�U�R����P�M��Bh��;��A����E�E��  �E�_^[���   ;��%�����]� ���������������������������������������������������������U����   SVW��@����0   ������j h�  h0��M�K����0�_^[���   ;�������]����������������������U����   SVW��@����0   ������j h�  h0��M������0�_^[���   ;��?�����]����������������������U����   SVW��@����0   ������h� �M�T�����tj h�  h0��M�Z������s����h��h0�貽�����0�_^[���   ;�������]������������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B��;��B���_^[���   ;��2�����]� ����������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bx��;������_^[���   ;��������]������������������������������U����   SVW��(����6   ������j h�  h0���,���P�M芳�����������,���蹳���0�_^[���   ;��F�����]�����������������������������U����   SVW��(����6   ������j h�  h0���,���P�M�
������}�����,����9����0�_^[���   ;��������]�����������������������������U���  SVW�������B   ��������3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |I�E�M������E��E���
}�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�먋E��D� j �E�P�M�����ER��P� r�ɷ��XZ_^[�M�3��%�����  ;�������]�   (r����   4rhexstring ����������������������������������������������������������������������������������U���  SVW��x����b   ������} ��   �}   @��   j h�������������Pj0j jj �E�U�観����x�����|���߭x����5�����$������P�ڴ����P�MQ���������������������������E�^  �  �} ��   �}   ��   j h���������(���Pj0j jj �E�U�
������x�����|���߭x����5�����$������P�<�����P�MQ�������������R����������G����E��   �r�} |l	�}   vaj h������������Pj0j jj �m�5�����$������P�ų����P�MQ�������������ۯ���������Я���E�Lj h��������4���P�EP��,���Q�z�����P�UR�V�������,���药�������肯���E_^[�Ĉ  ;�������]��������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   ��������E P�MQ�UR�EP���E�$��,���Q����B�H$�у�;�����P�M�e�����,����g����E_^[���   ;��������]���������������������������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ�������_^[���   ;��u�����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�f������E��}� u3��5�M������E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;�������]������������������������������������������U����   SVWQ��(����6   ������Y�M�j�v   ���E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;������_^[���   ;��������]� ���������������������������������������U����   SVW��@����0   ������h���EPh^� �������_^[���   ;��r�����]�������������������������U����   SVWQ��(����6   ������Y�M�j�v������E�}� t	�E�x u3����E�P�M�Q�҃�;������_^[���   ;��������]����������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u���� ��EP�MQ�U�R�E�H�у�;��b���_^[���   ;��R�����]� ��������������������������������������U���h  SVWQ��������   ������Y�M�j�F������E�}� t	�E�x u�M�w����E�2��EP�M�Q������R�E�H�у�;������b   ���}�E_^[��h  ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������M���`�����M����   �����M���   �����E���ݘ�  �E�_^[���   ;��������]���������������������������������������������U���L  SVWQ�������S   ������Y�M��M��R����M����G����M���0�<����M���H�1��������$�����$�����$�����������M����P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������軴���M������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������p����M���0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������%����M���H���P�Q�P�Q�P�Q�P�Q�@�A�E�_^[��L  ;��>�����]�����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E����X�M����Y�U�����E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��E��E��E�X�E��E�X�E�_^[��]� �����������������������U����   SVWQ��(����6   ������Y�M�j�6������E�}� t	�E�x u� ��EP�MQ�U�R�E�H�у�;�赽��_^[���   ;�襽����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u�$��EP�MQ�UR�E�P�M�Q�҃�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��(����6   ������Y�M�j ��������E�}� t	�E�x  u3��$��EP�MQ�UR�E�P�M�Q �҃�;��o���_^[���   ;��_�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j$�V������E�}� t	�E�x$ u3����EP�M�Q�U�B$�Ѓ�;��׻��_^[���   ;��ǻ����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x( u�(��EP�MQ�UR�EP�M�Q�U�B(�Ѓ�;��-���_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u��� ��EP�MQ�U�R�E�H,�у�;�蓺��_^[���   ;�胺����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j0�v������E�}� t	�E�x0 u3��)����E�$�EP�MQ�U�R�E�H0�у�;�����_^[���   ;��ڹ����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4��������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��K���_^[���   ;��;�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8�6������E�}� t	�E�x8 u���E�P�M�Q8�҃�;�轸��_^[���   ;�譸����]������������������������������������U���@  SVWQ�������P   ������Y�M�jD�������E�}� t	�E�xD u�M�ͻ���E�.��E�P������Q�U�BD�Ѓ�;������   ���}�E_^[��@  ;��������]� ������������������������������������������������U����   SVWQ��(����6   ������Y�M�jH��������E�}� t	�E�xH u���EP�M�Q�U�BH�Ѓ�;��i���_^[���   ;��Y�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jL�V������E�}� t	�E�xL u������EP�M�Q�U�BL�Ѓ�;��ֶ��_^[���   ;��ƶ����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�jP�������E�}� t	�E�xP u���EP�M�Q�U�BP�Ѓ�;��9���_^[���   ;��)�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jT�&������E�}� t	�E�xT u���EP�M�Q�U�BT�Ѓ�;�詵��_^[���   ;�虵����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jX�������E�}� t	�E�xX u3��4��E P�MQ�UR�EP�MQ�UR�EP�M�Q�U�BX�Ѓ� ;������_^[���   ;�������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j`��������E�}� t	�E�x` u3����E�P�M�Q`�҃�;��k���_^[���   ;��[�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jd�V������E�}� t	�E�xd u3����EP�M�Q�U�Bd�Ѓ�;��׳��_^[���   ;��ǳ����]� �������������������������������������������U����   SVWQ������:   ������Y�M�jh�������E�}� t	�E�xh u�M�����E�:��EP�M�Q�����R�E�Hh�у�;��'���P�M���������艰���E_^[���   ;�� �����]� ����������������������������������������������������U����   SVWQ��(����6   ������Y�M�jp��������E�}� t	�E�xp u������E�P�M�Qp�҃�;��j���_^[���   ;��Z�����]���������������������������������U����   SVWQ��(����6   ������Y�M�jl�V������E�}� t	�E�xl u������E�P�M�Ql�҃�;��ڱ��_^[���   ;��ʱ����]���������������������������������U����   SVWQ��(����6   ������Y�M�jt��������E�}� t	�E�xt u3����E�P�M�Qt�҃�;��K���_^[���   ;��;�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jx�6������E�}� t	�E�xx u���EP�M�Q�U�Bx�Ѓ�;�蹰��_^[���   ;�詰����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j|�������E�}� t	�E�x| u���E�P�M�Q|�҃�;��-���_^[���   ;�������]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u���E�P�M싑�   �҃�;�蔯��_^[���   ;�脯����]�������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u������EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;��ݮ����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��J���_^[���   ;��:�����]� ����������������������������������������������U����   SVWQ������<   ������Y�M�h�   �#������E�}� t�E샸�    u�M�c����E�9��E�P�����Q�U싂�   �Ѓ�;�蒭��P�M�ڶ��������ܕ���E_^[���   ;��k�����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u������E�P�M싑�   �҃�;��Ѭ��_^[���   ;��������]����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u���EP�M�Q�U싂�   �Ѓ�;��0���_^[���   ;�� �����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;�膫��_^[���   ;��v�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��ڪ��_^[���   ;��ʪ����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��2���_^[���   ;��"�����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��+��EP�MQ�UR�EP�M�Q�U싂�   �Ѓ�;�肩��_^[���   ;��r�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u����#��EP�MQ�U�R�E싈�   �у�;��٨��_^[���   ;��ɨ����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��*���_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��v���_^[���   ;��f�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��Ʀ��_^[���   ;�趦����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u������EP�M�Q�U싂�   �Ѓ�;�����_^[���   ;�������]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;�肥��_^[���   ;��r�����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����E�P�M싑�   �҃�;�����_^[���   ;��Ҥ����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��B���_^[���   ;��2�����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����E�P�M싑�   �҃�;�袣��_^[���   ;�蒣����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��'��EP�MQ�UR�E�P�M싑�   �҃�;������_^[���   ;�������]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��R���_^[���   ;��B�����]�����������������������������������������U����   SVWQ������>   ������Y�M�h�   �3������E�}� t�E샸�    u�M耤���E�N��EP�M�Q�����R�E싈�   �у�;�螡���U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��f�����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u�#��EP�MQ�U�R�E싈�   �у�;�輠��_^[���   ;�謠����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�P�M싑�   �҃�;��"���_^[���   ;�������]�����������������������������������������U����   SVWQ������>   ������Y�M�h�   �������E�}� t�E샸�    u�M�P����E�N��EP�M�Q�����R�E싈�   �у�;��n����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��6�����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u�#��EP�MQ�U�R�E싈�   �у�;�茞��_^[���   ;��|�����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����E�P�M싑�   �҃�;�����_^[���   ;�������]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��N���_^[���   ;��>�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u���#��EP�MQ�U�R�E싈�   �у�;�誜��_^[���   ;�蚜����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u�,����E�$�EP�MQ�U�R�E싈�   �у�;�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�U�R�E싈�   �у�;��J���_^[���   ;��:�����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;�螚��_^[���   ;�莚����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h   �������E�}� t�E샸    u3����EP�M�Q�U싂   �Ѓ�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h  ��������E�}� t�E샸   u3����E�P�M싑  �҃�;��b���_^[���   ;��R�����]�����������������������������������������U����   SVWQ������>   ������Y�M�h  �C������E�}� t�E샸   u�����$�M蕎���E�J��E�P�����Q�U싂  �Ѓ�;�誘���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��r�����]� ������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��E�X�M��E�Y�U��E��E�_^[��]� �����������������������U����   SVWQ������>   ������Y�M�h  ��������E�}� t�E샸   u�����$�M�E����E�J��E�P�����Q�U싂  �Ѓ�;��Z����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��"�����]� ������������������������������������������������������U����   SVWQ������>   ������Y�M�h  �������E�}� t�E샸   u�����$�M�U����E�J��E�P�����Q�U싂  �Ѓ�;��j����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��2�����]� ������������������������������������������������������U����   SVWQ��(����6   ������Y�M�h  �������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;�萕��_^[���   ;�耕����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h  �s������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;�����_^[���   ;��������]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h  ��������E�}� t�E샸   u���EP�M�Q�U싂  �Ѓ�;��P���_^[���   ;��@�����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�h   �3������E�}� t�E샸    u3����E�P�M싑   �҃�;�貓��_^[���   ;�袓����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h$  �������E�}� t�E샸$   u3����EP�M�Q�U싂$  �Ѓ�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h(  ��������E�}� t�E샸(   u3��'��EP�MQ�UR�E�P�M싑(  �҃�;��f���_^[���   ;��V�����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h,  �C������E�}� t�E샸,   u�'��EP�MQ�UR�E�P�M싑,  �҃�;�踑��_^[���   ;�訑����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h0  �������E�}� t�E샸0   u3����E�P�M싑0  �҃�;�����_^[���   ;�������]�����������������������������������������U����   SVWQ��(����6   ������Y�M�h4  ��������E�}� t�E샸4   u3����EP�M�Q�U싂4  �Ѓ�;��n���_^[���   ;��^�����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h8  �S������E�}� t�E샸8   u3��#��EP�MQ�U�R�E싈8  �у�;��ʏ��_^[���   ;�躏����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h<  �������E�}� t�E샸<   u�'��EP�MQ�UR�E�P�M싑<  �҃�;�����_^[���   ;�������]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h@  ��������E�}� t�E샸@   u�'��EP�MQ�UR�E�P�M싑@  �҃�;��h���_^[���   ;��X�����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�hD  �C������E�}� t�E샸D   u3����E�P�M싑D  �҃�;����_^[���   ;�貍����]�����������������������������������������U����   SVWQ��(����6   ������Y�M�hH  �������E�}� t�E샸H   u3����EP�M�Q�U싂H  �Ѓ�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�hL  �������E�}� t�E샸L   u3��#��EP�MQ�U�R�E싈L  �у�;��z���_^[���   ;��j�����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�hP  �S������E�}� t�E샸P   u3��'��EP�MQ�UR�E�P�M싑P  �҃�;��Ƌ��_^[���   ;�趋����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�hT  �������E�}� t�E샸T   u���'��EP�MQ�UR�E�P�M싑T  �҃�;�����_^[���   ;�������]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�hX  ��������E�}� t�E샸X   u�0����E�$�EP�MQ�UR�E�P�M싑X  �҃�;��_���_^[���   ;��O�����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j<�F������E�}� t	�E�x< u� ��EP�MQ�U�R�E�H<�у�;��ŉ��_^[���   ;�赉����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M�j@�������E�}� t	�E�x@ u3����EP�M�Q�U�B@�Ѓ�;��'���_^[���   ;�������]� �������������������������������������������U����   SVW��4����3   ������j�K   ���E��}� u3���E���H��;�蠈��_^[���   ;�萈����]�����������������������U����   SVW��@����0   ������h���EPh�� 耘����_^[���   ;��2�����]�������������������������U����   SVW��(����6   ������E�8 u�>j�q������E��}� u�)�E��M��E�P�M��Q�҃�;�蹇���E�     R��P�<��u��XZ_^[���   ;�菇����]Ð   D�����   P�i ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3��$��EP�MQ�UR�EP�U�M��B��;��߆��_^[���   ;��φ����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u���EP�MQ�U�M��B��;��I���_^[���   ;��9�����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j�v������E�}� t	�E�x u���EP�MQ�U�M��B��;�蹅��_^[���   ;�詅����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3��,��EP�MQ�UR�EP�MQ�UR�E�M��P��;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �6������E�}� t	�E�x  u3��(��EP�MQ�UR�EP�MQ�U�M��B ��;��k���_^[���   ;��[�����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u3��$��EP�MQ�UR�EP�U�M��B$��;�迃��_^[���   ;�诃����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3��$��EP�MQ�UR�EP�U�M��B(��;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�F������E�}� t	�E�x, u3��6��E$P���E�$���E�$�MQ�UR�EP�U�M��B,��;��m���_^[���   ;��]�����]�  �������������������������������������������������U����   SVWQ��(����6   ������Y�M�j0�������E�}� t	�E�x0 u3��(��EP�MQ�UR�EP�MQ�U�M��B0��;�軁��_^[���   ;�諁����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4��������E�}� t	�E�x4 u3��9��E(P���E �$�MQ�UR�EP�MQ�UR�EP�U�M��B4��;������_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u�����EP�MQ�U�M��B8��;��W���_^[���   ;��G�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�v������E�}� t	�E�x< u���EP�MQ�U�M��B<��;����_^[���   ;������]� �����������������������������U����   SVWQ��(����6   ������Y�M�j@��������E�}� t	�E�x@ u3����EP�MQ�U�M��B@��;��'��_^[���   ;������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jH�F������E�}� t	�E�xH u3����EP�MQ�U�M��BH��;��~��_^[���   ;��w~����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jD�������E�}� t	�E�xD u3����EP�MQ�U�M��BD��;���}��_^[���   ;���}����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jL�������E�}� t	�E�xL u���!��EP���E�$�U�M��BL��;��B}��_^[���   ;��2}����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jP�f������E�}� t	�E�xP u3����EP�MQ�U�M��BP��;��|��_^[���   ;��|����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jT��������E�}� t	�E�xT u3��$��EP�MQ�UR�EP�U�M��BT��;���{��_^[���   ;���{����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�jX�&������E�}� t	�E�xX u3��,��EP�MQ�UR�EP�MQ�UR�E�M��PX��;��W{��_^[���   ;��G{����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u3��,��EP�MQ�UR�EP�MQ�UR�E�M��P\��;��z��_^[���   ;��z����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u蒆���M��A�E��x u3���E�P�MQ�UR�EP�M��I��i��_^[���   ;���y����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�EP�MQ�U��J��o���E���P��y����_^[���   ;��hy����]� ����������������������������U����   SVWQ��4����3   ������Y�M��E��x u�r����M��A�E��x t�EP�MQ�U��J��^��_^[���   ;���x����]� ���������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t+�MQ�UR�EP�MQ�UR�EP�M��I�(�����0����
ǅ0���    ��0���_^[���   ;��?x����]� �����������������������������������U����   SVWQ��0����4   ������Y�M��E��x t'�MQ�UR�EP�MQ�UR�E��H�6�����0����
ǅ0���    ��0���_^[���   ;��w����]� ���������������������������������������U����   SVWQ��0����4   ������Y�M��E��x u袃���M��A�EP�MQ�UR�EP�M��k����u3��<�E��x t#�MQ�UR�EP�MQ�U��J��u����0����
ǅ0���    ��0���_^[���   ;���v����]� �������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t#�MQ�UR�EP�MQ�U��J�[t����0����
ǅ0���    ��0���_^[���   ;��'v����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t5�M$Q���E�$���E�$�UR�EP�MQ�U��J�|i����0����
ǅ0���    ��0���_^[���   ;��uu����]�  �����������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t'�MQ�UR�EP�MQ�UR�E��H��q����0����
ǅ0���    ��0���_^[���   ;���t����]� ���������������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;��gt��_^[���   ;��Wt����]������������������������������U����   SVW��@����0   �������EP����Q��P  �Ѓ�;���s��_^[���   ;���s����]������������������������������U����   SVW��(����6   ������} u3��m�EP�ev�����E��}� u3��T��E��M��I �PP��;��ns���E�}� uh�������P�x\����3����E�M�I ���   ��;��1s��_^[���   ;��!s����]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;��mr��_^[���   ;��]r����]��������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;��r��_^[���   ;���q����]��������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;��mq���M��A�E����M��   _^[���   ;��Gq����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;���p���M��A�E����M��   _^[���   ;���p����]� ���������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ������9   ������Y�M��E�E�}� t�E��U�<� u3��W�E����M��B��;��Oo��P�M�:����E���j �E��U��P�M�Q�U���M��P��;��o����u3���   _^[���   ;���n����]� ��������������������������������������������������U����   SVWQ������<   ������Y�M��E�E�}� t�E��U�<� u3��G�E��U��P�M����M��B��;��cn��P������}z��P�M��T���������w���   _^[���   ;��.n����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�MQ�U�R������   �Q\�҃�;��m���E�_^[���   ;��m����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M�j �E�P�M�x���E�_^[���   ;��m����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�UR������   �Q�҃�;��l��_^[���   ;��l����]� �������������������������������U����   SVWQ������9   ������Y�M��E��x�u3��   �E��x t�E��@�   �E�    j�g�����E���M��u���E��}� t8�M��(]���E�E����M��B��;���k���M�9u�E��M�H�E��$�h�������P��T�����E��@����3�_^[���   ;��k����]���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B(��;��k��_^[���   ;��k����]������������������������������U����   SVWQ������9   ������Y�M��E����M��B��;��j��9Eu�} u�   �<�EP�MQ�� ����v��P�M�Q���� ����t���M�m����t3���   _^[���   ;��Oj����]� ���������������������������������������������������U����   SVWQ��4����3   ������Y�M�j�E�Q�S���������_^[���   ;���i����]� ���������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M�j�E�Q�Ma���������_^[���   ;��i����]� ���������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M�j�E�Q�8M���������_^[���   ;��mh����]� ���������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U���  SVW��������   ������} u3��  �E���M�B��;��g���E�j h@  ������P�Ek�����E�������E������ǅ�����?�E������ǅ����l6ǅ�����5ǅ����7*ǅ ���)ǅ����Aǅ����9ǅ���U*ǅ���%ǅ����5ǅ����9ǅ���)ǅ ����/ǅ$���#%ǅ(���))ǅ,���)ǅ0����/ǅ4���S,ǅ8����/ǅ<����/ǅ@����,ǅD���R(ǅH����)ǅL���d%ǅP���%ǅT���<*ǅX���%ǅ\���i%h@  ������P�MQ�U�Rj�w_����R��P�P��S��XZ_^[��  ;��ze����]�   X�����@  d�np �������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��JN���E�� L��E��M�H�E��M�H�E�_^[���   ;��d����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M���J���E��t�E�P�iR�����E�_^[���   ;��d����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���V��_^[���   ;��c����]������������������U����   SVWQ��4����3   ������Y�M��E��P�E��H��I �R`��;��fc��_^[���   ;��Vc����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��P�E��H��I �R\��;���b��_^[���   ;���b����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�M��Q�E��H�I �Rd��;��b��_^[���   ;��rb����]� ����������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U��B�M��Q�J ���   ��;��a��_^[���   ;��oa����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�M��Q�J ���   ��;���`��_^[���   ;���`����]� �������������������������������U���  SVW��l����e   ������} u3��   �E���M�B��;��`���E�j h�   ��0���P��d�����E��P����E��0���ǅ4����?�E��p���ǅt����5ǅx���7*ǅ|���l6�E��,�E�)�E��Ah�   ��0���P�MQ�U�Rj��Y����R��P�����M��XZ_^[�Ĕ  ;���_����]ÍI     �0����   �np ��������������������������������������������������������������������������������̋�`<����������̋�`L����������̋�`l����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`P����������̋�``����������̋�`p����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`d����������̋�`t����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`X����������̋�`h����������̋�`����������̋�`����������̋�`,�����������U����   SVW��@����0   ���������H���   ��;��]��_^[���   ;��o]����]����������������������U����   SVW��@����0   �������E�Q����B���   �у�;��]���E�     _^[���   ;���\����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q���   �Ѓ�;��\��_^[���   ;��\����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B���   �у�;��\��_^[���   ;��\����]� ����������������������������������U����   SVW��@����0   ���������H����;��[��_^[���   ;��[����]��������������������������U����   SVW��@����0   �������E�Q����B�H�у�;��H[���E�     _^[���   ;��/[����]��������������������������������������U����   SVW��@����0   �������E�Q����B�H�у�;���Z���E�     _^[���   ;��Z����]��������������������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q����B���   �у�;��6Z������g��������� ����c�������_^[���   ;��Z����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��Y��_^[���   ;��Y����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H\�у�;��!Y��_^[���   ;��Y����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H���   �҃�;��X��_^[���   ;��X����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�HX�у�;��X��_^[���   ;���W����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B �Ѓ�;��W��_^[���   ;��W����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B���   �у�;��W��_^[���   ;��W����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;��V��_^[���   ;��yV����]� �����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��   �у�;��V��_^[���   ;���U����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��B$��;��U��_^[���   ;��yU����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H(�у�;��U��_^[���   ;���T����]� �������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q�B`�Ѓ�(;��qT��_^[���   ;��aT����]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H,�у�;���S��_^[���   ;���S����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��^����P�M���a����Pj j �E�P����Q�B4�Ѓ� ;��MS��_^[���   ;��=S����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���R��_^[���   ;���R����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��eR��_^[���   ;��UR����]����������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H4�у� ;���Q��_^[���   ;���Q����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q@�҃�;��^Q��_^[���   ;��NQ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HD�у�;���P��_^[���   ;���P����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;��eP��_^[���   ;��UP����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;���O��_^[���   ;���O����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BP�Ѓ�;��O��_^[���   ;��uO����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;��O��_^[���   ;��O����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;��N��_^[���   ;��N����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���   �҃�;��N��_^[���   ;���M����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P����Q���   �Ѓ�;��M��P�M��M���� �����V���E_^[���   ;��\M����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�Bh�Ѓ�;���L��_^[���   ;���L����]����������������������������U����   SVW��0����4   ������hx������Ph��h�   �)T������8�����8��� t��8����Y����0����
ǅ0���    ��0���_^[���   ;��FL����]���������������������������������������������U����   SVW��$����7   ������E�8 t?�E���8�����8�����,�����,��� tj��,�����V����$����
ǅ$���    �E�     _^[���   ;��K����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��M���<���E��t�E�P�i9�����E�_^[���   ;��K����]� ������������������������U����   SVWQ��4����3   ������Y�M��M����oD���M��/O���E�_^[���   ;��J����]��������������������U����   SVWQ��(����6   ������Y�M��M���Q���E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��0J����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M���B���M�����?��_^[���   ;���I����]�����������������������U����   SVWQ��4����3   ������Y�M��M��9��_^[���   ;��kI����]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E����Xp�E��@x�����E��@|   _^[��]������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	�2O���E��     �E��x` t�E���`P�1����_^[���   ;��SH����]������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 thx������P�1�����E��x` thx������P��0�����M���@���M��%L���E�P�M���dQ�U��BxP�MQ�U���`R�rP�����M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�f0�����E��@|�   �E��xd ��   �E���pP�M���hQ�UR�BE������u(�E��@h    �E����Xphx������P�0�����EP�M����P��j j j�E���P�M��	�qM���U��B|�E��x|t�M��?���E��@|��E��@x�����E��@|_^[���   ;��F����]� ������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M���>���M��BJ��_^[���   ;���E����]��������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	��K���U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;���D����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap��E��xd t�E��@h��E��x|u�   �3�_^[��]� ��������������������������������U����   SVW��@����0   ���������H����;���C��_^[���   ;���C����]��������������������������U����   SVW��@����0   �������E�Q����B�H�у�;��C���E�     _^[���   ;��oC����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H�у� ;���B��_^[���   ;���B����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;��qB��_^[���   ;��aB����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���A��_^[���   ;���A����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q�҃�;��~A��_^[���   ;��nA����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M���'�����M��'���H �G@��;���@��_^[���   ;���@����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��2'�����M��('���H �GD��;��d@��_^[���   ;��T@����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M��&���xH u3��#�M��&�����M��&�����H �FH��;���?��_^[���   ;��?����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M�� &���xL u3��/��EP�MQ�UR�M�� &�����M���%���H �GL��;��2?��_^[���   ;��"?����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M��%���xP u����3��EP�MQ�UR�EP�M��[%�����M��Q%���H �WP��;��>��_^[���   ;��}>����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M���$���xT u����+��EP�MQ�M���$�����M��$���H �WT��;���=��_^[���   ;���=����]� �����������������������������������������U���  SVWQ�������C   ������Y�M��} t<�M��5$����E�P�M��,$�����M��"$���H �WL��;��^=���M��M���&���} t?��������B��P�M�n)���������%���M���#���@@�EЃ}� t�E�P�M�C)��R��P���� +��XZ_^[��  ;���<����]� �I    ������   ��bc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��#���x` u� }  �'��EP�M���"�����M���"���H �W`��;��'<��_^[���   ;��<����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��j"�����M��`"���H �WH��;��;��_^[���   ;��;����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�j�EP��E���������P�M��Y&���E�M�I��;E��M�+F��;E�~������3��EP�MQ�UR�EP�M��!�����M��!���H �WD��;���:��_^[���   ;��:����]� ���������������������������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M��� ���xP u������;��EP�MQ�UR�EP�MQ�UR�M�� �����M�� ���H �GP��;���9��_^[���   ;���9����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��  ���xT u������+��EP�MQ�M�� �����M������H �WT��;��39��_^[���   ;��#9����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M�����xX u�'��EP�M��j�����M��`���H �WX��;��8��_^[���   ;��8����]� ��������������������������������U����   SVW�� ����8   ������M��?4���E�P�MQ�5E������t�}� u3���E�P�M�Q�U�R�E�P�M��L<��R��P����%��XZ_^[���   ;���7����]ÍI    �����   �dat ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVWQ������<   ������Y�M��M�^���M���+����uhx������P������3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;��~6����u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�l���͍E�P��-�����   R��P���$��XZ_^[���   ;��6����]�    �����   �����   �arr count ����������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M��!���M��T*����uhx������P�b����3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;���4����u3��i�}� u3��_�E�    �	�Eԃ��EԋE�;E�}4�EԋM��<� t�EԋM����)����u�ϋEԋM���R�M�<��뻍E�P�C,�����   R��P�`�"��XZ_^[���   ;��l4����]�    h����   �����   �arr count ��������������������������������������������������������������������������������������U����   SVW��@����0   ���������H��   ��;��3��_^[���   ;��3����]����������������������U����   SVW��@����0   �������E�Q����B��$  �у�;��E3���E�     _^[���   ;��,3����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��(  �у�;��2���E�_^[���   ;��2����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��,  �у�;��>2��_^[���   ;��.2����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��,  �у�;��1�������_^[���   ;��1����]� ���������������������������U����   SVW��@����0   ���������H��0  ��;��O1��_^[���   ;��?1����]����������������������U����   SVW��@����0   ���������H��4  ��;���0��_^[���   ;���0����]����������������������U����   SVWQ��0����4   ������Y�M��} t�M�5,����0����
ǅ0���    ��0���P�M�Q����B��8  �у�;��[0��_^[���   ;��K0����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��<  �у�;���/��_^[���   ;��/����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q��@  �Ѓ�;��F/��_^[���   ;��6/����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H��D  �҃�;���.��_^[���   ;��.����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��H  �у�;��N.��_^[���   ;��>.����]� ����������������������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R����H��L  �҃�;���-��P�M�7���� �������E_^[���   ;��-����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��T  �Ѓ�;��2-��_^[���   ;��"-����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��P  �Ѓ�;���,��_^[���   ;��,����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��X  �у�;��N,��_^[���   ;��>,����]� ����������������������������������U����   SVW��@����0   ���������H��\  ��;���+��_^[���   ;���+����]����������������������U����   SVW��@����0   �������E�Q����B��`  �у�;��u+���E�     _^[���   ;��\+����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��d  �҃�;���*��_^[���   ;���*����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��h  �҃�;��O*��_^[���   ;��?*����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M����_^[���   ;���)����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��{)����]������������������U����   SVWQ��4����3   ������Y�M��EP�M��
��_^[���   ;��')����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M��7��_^[���   ;���(����]������������������U����   SVWQ��4����3   ������Y�M�jh�  �M�$���EP�MQ�M���!��_^[���   ;��d(����]� ������������������������U����   SVWQ��(����6   ������Y�M��E����M��BX��;��(��P�M�O����t$ǅ,���   ��,���P�MQ������   ��EP�MQ�UR�EP�M���!��_^[���   ;��'����]� ����������������������������������������U����   SVWQ��0����4   ������Y�M�j �M�	'��� ��0�����0����  t�7�5�3�E��x u*j h�  �M�W$����uj h�  �M�D$����t3�� �EP�MQ�UR�EP�MQ�UR�M��#,��_^[���   ;���&����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��^&��_^[���   ;��N&����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �EP�����_^[���   ;���%����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��@   �   _^[��]� ���������������������U����   SVWQ��4����3   ������Y�M��E��@   _^[��]� ��������������������������U���`  SVWQ�������X   ������Y�M��}`��u
�E��@   �}��   �E�E�j �M��v$���8�  u)�2��P�M��	&��jh�  �M�2 ���   �  �vj �M��;$���8�  u*��EP�MQ�U���M��P��;��e$���   �j  �:j �M���#���8�  tj �M���#���8ujh�  �M����E��@    �}�  �E�E��E��H���U��Jj	�E����M��BX��;���#��P�a1�����E��E�    �}� tj �M��(���EȋE��M�;H��  �E��x ��  j h�  �M�� ����uj h�  �M� �����s  j h�  �M�����}� tj �M��D(���EȋE��MȉH�M��(���} t�M������uǅ����   �M��}���������)  �EP� �����M�����j�M�����P�M�����t�������E��|����M�����E��E��t����E�   �M�-��������������t������t������t��E�   ��E�   ��E�   ��E�    ������t��� t��t��������t���P�M����M��BX��;��A"��P�������t��� t��t����N����t����U'���M��M'���M��a���EP�MQ�UR�EP�M��#��R��P������XZ_^[��`  ;���!����]�    ����   .����   +t���   (md mu pActive ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��^ ��_^[���   ;��N ����]� ����������������������������������U����   SVW��4����3   ������j�   ���E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;����_^[���   ;������]����������������������������������������������U����   SVW��@����0   ������h���EPh�f �/����_^[���   ;��2����]�������������������������U����   SVW������<   ������j�{������E��}� t	�E��x uǅ��������M�]��������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�_(���EP�M��Q�҃�4�� ����M����� ���_^[���   ;��m����]����������������������������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;�����_^[���   ;�������]�����������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�M��Q�҃�;��P��_^[���   ;��@����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� ���M��>��_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M��M��A���E��t�E�P�
�����E�_^[���   ;��d����]� ������������������������U����   SVWQ��(����6   ������Y�M��M�w���E�M��Q�P�E�M��Q�P�E�    �	�E���E�E��M�;H}�E��H�U��P�M�����u3���͸   _^[���   ;������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��} |$�E��M;H}�} |�E��M;H}�E;Eu�"�E��H�U��P�M��Q�E��Q�z����_^[���   ;������]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E;E}	�E���E�} |$�E��M;H}�} |�E��M;H}�E;Eu�/�E��H�U���E�EP�M������t�EP�M�Q�M����_^[���   ;��7����]� �������������������������������������������U����   SVWQ������9   ������Y�M��E��x u�E��H�M��%�E��x t�E��H�U�J�M���E��H��M��}� u3��]��h������P�M���Q�U��BP����Q��  �Ѓ�;��g���E�}� u3���E��M�H�E��M��H�   _^[���   ;��3����]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��P;Qu�M������u3��&�E��H�U��B�U���E��H���U��J�   _^[���   ;������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��M;H}�EP�MQ�M�� ���#�E��H;M}j �M�������EP�M�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3���E��H�U�E���   _^[��]� ���������������������������U����   SVWQ��(����6   ������Y�M��E��M;H~	�E��H�M�} }�E    �E��M��P;Qu�M������u3��Z�E��H�M��	�E���E�E�;E~�E��H�U��B�U�u�L�����ԋE��H�U�E���E��H���U��J�   _^[���   ;��z����]� ��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3��E�E��H���U��J�	�E���E�E��M;H}�E��H�U��B�U�u�L����Ѹ   _^[��]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M����P�M����_^[���   ;��>����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E��M�;H}�E��H�U��;Eu�E���ԃ��_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E���P������E��@    �E��@    �M��A    _^[���   ;��6����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��@    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M��E��H��Q�M���#���E�}� t�E��H��Q�M������E�_^[���   ;��c����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H}�E��H�U���3�_^[��]� �������������������U����   SVWQ��$����7   ������Y�M��EP�M���!��j�E��HQ�U��BP�M��K���R��P�P)� ��XZ_^[���   ;��~����]� ��   X)����   d)sort ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��4����E�� 4��E��M�H�E�_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�Ѓ�;����_^[���   ;��w����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�� @��E�_^[��]���������������������������U����   SVWQ��$����7   ������Y�M��EP�M��	 ��j�E��HQ�U��BP�MQ�M����R��P�4+����XZ_^[���   ;������]� ��   <+����   H+sort �����������������������������������U����   SVWQ��4����3   ������Y�M��E�� L��M�������M�������E��@    �M������E�_^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M��E�� X��E��@    �E��@    �E�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��M�����E��t�E�P�i������E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P��������E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� L��M��[���M�������M������_^[���   ;��,����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E����M��A�E����M��A�E��@    _^[��]���������������������������U���   SVWQ�� ����@   ������Y�M��M�����E��}� tm�M�����E�}� tM�E��������������������� t%��j��������������;������ ����
ǅ ���    �E�    �E�E�덋M������_^[��   ;�������]����������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t�M��Q�z t�E��H��0����
ǅ0���    ��0���_^[��]������������������������������������U����   SVWQ��0����4   ������Y�M��E����M�9At�U��B��0����
ǅ0���    ��0���_^[��]���������������������������U����   SVWQ������9   ������Y�M��M�����E��}� t�M��!���E�M�����E�E���_^[���   ;��W����]������������������������������U����   SVWQ������:   ������Y�M��E�    �M��$���E��}� tD�E�M�U���U�;�uǅ���   �
ǅ���    ����� t�E���M��c���E��3�_^[���   ;��
����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E�M��Q�P�E����M�A�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E����M�A�E�M��Q�P�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ������9   ������Y�M��E�    �M��d���E���M������E��}� t�E���E���E�_^[���   ;��	����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� X��M�����_^[���   ;������]�������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E�H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t;�E��x t2�E��H�U��B�A�E��H�U��B�A�E��@    �M��A    _^[��]�����������������������������������U����   SVW��4����3   ������E��M��E�M���E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M����_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��M�%���E_^[���   ;��h����]� ����������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]�  ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��(����6   ������Y�M��} u3��]��EP�M���M��B@��;�����E�}� u3��6�M��J�����P�EP�MQ����B0���   �у�;�����M�����_^[���   ;��l����]� ������������������������������������������������U����   SVWQ������=   ������Y�M���EP����Q0�B�Ѓ�;������E�}� tM�E쉅 ����� ������������� t%��j��������������;����������
ǅ���    �E�    _^[���   ;������]� ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�j�E�Q���������t�   �3�_^[���   ;�� ����]� ��������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�j�E�Q���������t�   �3�_^[���   ;�� ����]� ��������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��c���_^[���   ;��S�����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;������_^[���   ;��������]����������������������������������U����  SVW��(����v   ������ǅ ���    �}( uǅ0���    �M�������0����!  �E�    �M��������  �M��B����M����������   �EP��H����G����� ���j h������������� ���P��l��������� ���j j���H���Q��l���R������P�E������� ���P������Q�q������� ���P������R�Z������� ��� P�M��������:�����uǅ(���   �
ǅ(���    ��(�����?����� ����� t�� ���ߍ������������ �����t�� �������������� �����t�� ���������������� �����t�� ������l��������� �����t�� �����������:����� �����t�� ������H����R�����?�����t(�E(P�M$Q�M��L���P�UR�EP�MQ�f������E��M��e���!�E(P�M$Qj �UR�EP�MQ�;������E��E�������M���������R��P��?�>���XZ_^[���  ;��)�����]ÍI    �?����   �?icon �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������EP�MQj �UR�EP�MQ�������_^[���   ;��
�����]���������������������������������U���  SVW��H����n   ������} u3��g  j h�   ��<���P���������$���P�M��M�B��;�������$��������t9j ��$���P�MQ�c�������u ǅL���    ��$���������L�����   �E��\����E��|����E�E��E��<���ǅ@����?�E��<�E��A�E�&@�E��-�E�=�E�A �E�� �E�!6�E��<�E��@�E�V=�E�0@�E�N@�E��<�E�R<�E�S@�Eĝ<�E�+@�E��A�E��-h�   ��<���P�MQ�URj	�G�������X�����$���������X���R��P��B�H���XZ_^[�ĸ  ;��3�����]Ð   �B<����   �B$���   �Bdescription np �������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B���   �у�;��2���_^[���   ;��"�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$���E�$�MQ�U�R����H���   �҃�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q���   �Ѓ�;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q���   �Ѓ�;��&���_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�Bp�Ѓ�;��5���_^[���   ;��%�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���  �҃�;��;���_^[���   ;��+�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���  �҃�;��;���_^[���   ;��+�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�� ����M���E�_^[���   ;��������]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P�������E��     _^[���   ;��^�����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]�����������������̋�`<����������̋�`L����������̋�`����������̋�` ����������̋�`0����������̋�`P����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`����������̋�`����������̋�`,�����������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M��f����E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��l�����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��<�����}�EP�M�Q�U�R�M��������U��������_^[��,  ;�������]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�������}�E�P�M�Q�U�R�M��3������U��������_^[��8  ;��n�����]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��#�����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��������}�E�P�M�Q�U�R�M��A������U��������_^[��8  ;�������]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��u�EP�MQ�UR�M������83��} ����t�EP�MQ�UR�M��������EP�MQ�UR�M�����_^[���   ;�������]� �������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  �Ek� E�E���E�P�MQ�U���M����;��{����Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;��
����Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��������t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;�������]� ����������������������������������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u�E� ����3���  �Ek� E�E���E�P�MQ�U���M����;������Eȃ}� u
�E��  ��}� }�E�     3��  �E�   �E���E��E�    �E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;��!����Eȃ}� uS�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��������t�
��E��E�뷋E���   ��}� }�Eԃ��E��	�Eԃ��E��D����}� ~�Eԃ��M���E�Mԉ�E�;M}F�E�M�M�M���E�P�MQ�U���M����;��U�����|h`������9P�d������E�8 ~I�E����MM�M���E�P�MQ�U���M����;�������h`������?P������3�_^[��  ;��������]� ������������������������������������������������������������������������������������������������������������������������������������������������������������u�U��� PRSVW�Ej P������_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR�R������E�@���E�;|�_^[��]���������������������������̋�U��V���t!��tS�]��tW�̋�����F�V�3_[^]� �������������̋�U��QSVW��3���;�tR�}�9>~K��    �F�8�����9T�u�D8�9t�N�T�ERP����������̋E�@���E�;|������̋u3��ƅ�tV�@G��u���tJ9u9Vu
9Vu9Vt�MWVQ����������̋F9T0�t�MWVQ����������̋vO��u�_^[��]� �����������������������������������������������������������̀=�� uj jj j j �������P�c�����������������������������jjj j j �s������������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������������̋�U��������} t������]�������̋�U�����10����*� ��F���:��7��10���J���F���(��[B]�������������������������������������̋�U��Q����E��M����E���]������������������̃=l ��������\$�D$%�  =�  u�<$f�$f��f���d$������ �~D$f(��f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�U������D$��~D$f��f(�f��=�  |!=2  �fT���\�f�L$�D$����f���fV��fT��f�\$�D$�������������������������������������������������������������������������������̃=` t-U�������$�,$�Ã=` t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������������������������������������������������������̋�U��Q�M��EP�M�Q��������]� ����������������̋�U��Q�M��E�� ��M�Q��������]��������������̋�U��Q�M��M������E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M�Q�M�������]� ����������������̋�U��Q�M��E�P���������]�������̋�U��Q�M��E���	P�M��	Q�|������������]� �������������������̋�U��Q�M��E���	P�M��	Q�<���������؋�]� ��������������������̋�U��Q�M��E���	P�M��	Q�������3҅���]� �����������������̋�U��Q�M��E�����]�������������̋�U��Q�M��E�� ��E���]� ��������������������̋�U��Q�M��E���]� �������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ����������������������������U��WV�u�M�}�����;�v;���  ���   r�=` tWV����;�^_u������   u������r)��$��b�Ǻ   ��r����$��a�$��b��$�Db��a b$b#ъ��F�G�F���G������r���$��b�I #ъ��F���G������r���$��b�#ъ���������r���$��b�I �b�b�b�b|btblbdb�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��b���b�b�b�b�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�Ld�����$��c�I �Ǻ   ��r��+��$�Pc�$�Ld�`c�c�c�F#шG��������r�����$�Ld�I �F#шG�F���G������r�����$�Ld��F#шG�F�G�F���G�������V�������$�Ld�I  dddd d(d0dCd�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�Ld��\dddtd�d�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋T$�L$��ti3��D$��u���   r�=` t�����W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̋�U��j�hx�h)d�    P���SVW���1E�3�P�E�d�    �}��   蝻����u3��  ������u�����3��  �������!����������������}���������3��i  �S�����|�������|j �`�������t�Q��������n���3��3  j���������������  �} um�=�� ~X���������E�    �=�� u�2���������/����	����E������   ��} u�=,��t������3��   �   �}��   �{���h�   h �jh  j�������E�}� tV�U�R�,�P�8�Q��!�Ѕ�t%j �U�R�H�������!�M��U��B�����j�E�P�;�����3���3����}u
j �8������   �M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��}u�����EP�MQ�UR�   ��]� �����������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �e��E�   �} u�=�� u3��N  �E�    �}t�}uT�=� t�EP�MQ�UR���E�}� t�EP�MQ�UR�S����E�}� u�E�    �E������E���   �EP�MQ�UR�"����E�}u=�}� u7�EPj �MQ�����URj �EP������=� t�MQj �UR���} t�}u@�EP�MQ�UR�������u�E�    �}� t�=� t�EP�MQ�UR���E��E������8�E���U��E�P�M�Q�������Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �����E�    �EP�Y   ���E��E������   �����ËE�M�d�    Y_^[��]������������������������������������������̋�U����TP��!�E��PQ��!�E��U�;U�r�E�+E�����s3���   j�M�Q�8������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}h\�j�E�P�M�Q�"������E��}� u:�U���U�E�;E�r%h�   h\�j�M�Q�U�R��������E��}� u3��Q�E�+E����M����U��E��E��M�Q��!�T�UR��!�M���U����U��E�P��!�P�E��]�����������������������������������������������������������������������������������������������̋�U��EP�����������؃�]��������������������̋�U��Qh�   h\�jjj ��������E��E�P��!�T�T�P�}� u�   ��U��    3���]�������������������������;��u��鯼������������������̋�U������]�h��  h?  �5������E��E%�  =�  ��   ���E�$�b������E�}�t�}�t!�}�t3�Jh��  �M�Q��������E�   h��  �U�R��������E���i�E�P���E�$j�}������P�M�Q�E������$���E�$jj�S������&�U������U�E�E�h��  �M�Q�_������E���]��������������������������������������������������������������������̺���A��������������������z�����������������̋�U��Qj j j���P�MQ�������E��E���]������������������������̋�U��j�EP�U�����]������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̋�U��Q�$�P��!�E��}� t�U�j�V�����jj �ʲ�����Z�����]�������������������̋�U��Q�E�    �$�P��!�E��MQ��!�$��E���]��������������̋�U��$�P��!]�������������̋�U��E��w$������4����tRP�EQP�D   ��]ú�R�   P�E�   QP�$   ��]�������������������������������̋�U���@  ���3ŉE��ES�]VW�}S������������ǅ����    �v�������������uS�������������5�!j j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ������h  ��  ����������t%��������L�PSQW�}  �����"  2��������� ������u���  ��t��!����   h  ������R������Ph  ������Q���S�:�������t-������������RWhH�������P�EQ������RP���   �=�!j j h
  ������Qj�������Rj h��  �0��ׅ�t������j j h
  ������Pj�������Qj h��  ���ׅ�t������������������������R�UPh��VQSR����������u̋M�_^3�[������]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@��!�	�   Ëe��E������E�M�d�    Y_^[��]��������������������������������������̋�U��j�h��h)d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@��!�	�   Ëe��E������E�M�d�    Y_^[��]����������������������������������������������������̋�U���  ���3ŉE��=����E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ��d�������A��u�Њ@��u�W������+�O�OG��u��������ȃ�����Ȋ@��u�������+���O�OG��u������ȃ��_������������SjPQ�������^[�M�3�������]��������������������������������������������������������������������̋�U���D  ���3ŉE�S���V�uW�}�����������   h��� "����   h��P��!������   ����   �M�Vh��QhL���$Rh@��~ Wh0�h��������h��Q�ЋV��$RW�E�P�M�Q��   ��8h���U�Rh���E�Ph��������Q��!������R��������������PjSQ������(_^[�M�3��G�����]�hP�jSW�������M�_^3�[�%�����]�����������������������������������������������������������������������������̋�U����ESV�u�E��EW3�+ƉE����M��r�   ;�s&�0�U���Qh��R���E��E����GF�ɋM�E�y� � _^[��]���������������������������������̋�U���  ���3ŉE��=����E��   SV����   �ȍq�A��u�+΃�:��   ww������3Ɋ���������A��u�Њ@��u�W������+�O�OG��u��������ȃ�����Ȋ@��u�������+���O�OG��u������ȃ��_�������SjP�EP������^[�M�3��_�����]�����������������������������������������������������������������������̸   ����������̋�U��E��w	����]�3�]������̋�U��M��w�U��������]Ã��]�����������̋�U��M������    ]�����������������̋�U��M������    ]�����������������̡�����������̡������������u�U��� PRSVWh0�h+�jBh��j蟬������u�_^[ZX��]������������������������̋�U���(]����̋�U���']����̋�U��j jh��h��h8�h   h   j �v�����P������]�������������������������̋�U��} u��EP�MQ�UR�EP�MQ�U���]������������������������̋�U��j �EP�K�����]�����������̋�U����EP�M��a����M�R�C�������et�E���E�M�R�ݩ������u�E�Q��������xu	�U���U�E��M��M�蕩������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M�������]������������������������������������������������̋�U��Q�M��E��@ �} ��   �"����M��A�U��B�M��Pl��E��H�U��Ah�B�M��;�t�E��H�Qp#H�u
�ɽ���M���U��B;H�t�M��Q�Bp#H�u�����M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������������������������������������������������������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]�������������������̋�U��Q�M��E���]����������������̋�U��j �EP�+�����]�����������̋�U���V�EP�M������M���t*�E�0�M��Y�������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��Ȧ������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M������^��]�������������������������������������������������������������������̋�U��Q�E�������Az	�E�   ��E�    �E���]���������������������̋�U����} t$�EP�MQ�U�R說�����E�M���U��P��EP�MQ�U�R�6������E�M���]������������������������������̋�U��j �EP�MQ�UR�������]�������������������̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�c�����3Ƀ} ���Mă}� u!h,�j h�  h��j蚥������u̃}� u3�M����    j h�  h��h��h,��M������   �  3�;E��ىM�u!hd�j h�  h��j�2�������u̃}� u3������    j h�  h��h��hd��������   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�������Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3�������]��������������������������������������������������������������������������������������������������������������������̋�U���@�E�    �E P�M��z���3Ƀ} ���M܃}� u!h,�j h3  h��j萣������u̃}� u@�C����    j h3  h��h��h,��C������E�   �M�������E���  3�;E��ىM�u!hd�j h4  h��j��������u̃}� u@������    j h4  h��h��hd��κ�����E�   �M��r����E��}  3��} ����#E��	;E��ىM�u!h(�j h<  h��j薢������u̃}� u@�I���� "   j h<  h��h��h(��I������E�"   �M�������E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�V  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��*�������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  h��h��hP�hH��U�R�E�P������P�8������M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE���X���t �U����0uj�M��Q�U�R跬�����E�    �M�������Eċ�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�B�����]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M�胬���} }�E    3Ƀ} ���M��}� u!h,�j h�  h��j茞������u̃}� u@�?����    j h�  h��h4�h,��?������E�   �M������E���  3�;E��ىM�u!hd�j h�  h��j��������u̃}� u@�ʽ���    j h�  h��h4�hd��ʵ�����E�   �M��n����E��g  �E�  �M��;M��ډU�u!h��j h�  h��j蘝������u̃}� u@�K���� "   j h�  h��h4�h���K������E�"   �M������E���  �M��Q�4�j���%�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ�������E��}� t�U� �E��E��M��b����E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ蕠�����E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M��ϼ���E���  �M��Q�?�J������� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4�һ��%�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M��B�������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U��֘���E�U��E܅���   �} ~}�M��Q���� #E�#U��M�莺��f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U��M����E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M�����f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4����%�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�ؘ������0�M��U���Uj h�  �E�P�M�Q�Q����E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q胘���Ѓ�0�E��M���Mj jd�U�R�E�P������E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�1����ȃ�0�U�
�E���Ej j
�M�Q�U�R譗���E��U��E���0�M��U���U�E�  �E�    �M������E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�Ӎ����]���������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�s�����3Ƀ} ���Mă}� u!h,�j h*  h��j誔������u̃}� u3�]����    j h*  h��hL�h,��]������   ��   3�;E��ىM�u!hd�j h+  h��j�B�������u̃}� u3������    j h+  h��hL�hd���������   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�A������Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�   ���EȋEȋM�3��Ӷ����]�����������������������������������������������������������������������������������������������������������̋�U���4�E�H���M��UR�M�襠��3��} ���E�}� u!h,�j h�  h��j軒������u̃}� u@�n����    j h�  h��hd�h,��n������E�   �M������E��  3�;U��؉E�u!hd�j h�  h��j�F�������u̃}� u@������    j h�  h��hd�hd���������E�   �M�蝲���E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P��  ���M��0�U����U���E�M�H�M��} ��   j�U�R�  ���M�蘐��� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�  ���EPj0�M�Q覑�����E�    �M��V����EЋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP蘯����]���������������̋�U���P���3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�?�����3Ƀ} ���M��}� u!h,�j ho  h��j�v�������u̃}� u3�)����    j ho  h��h|�h,��)������   �i  3�;E��ىM�u!hd�j hp  h��j��������u̃}� u3������    j hp  h��h|�hd���������   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�������E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�?������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ��������M�3�� �����]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ螭����]�����������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR輅�����E��{�}fu!�E P�MQ�UR�EP�MQ�7������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�-������E��#�U R�EP�MQ�UR�EP�MQ�۬�����E��E���]������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�����������������������̋�U��} t#�EP��������P�MQ�UUR������]����������������̋�U��Q�E�    �	�E����E��}�
s�M�����R��!�M������ԋ�]�����������������̋�U��} u� �    ��EP��!�x� �   ]��������������̋�U���`���3ŉE��E� �E� �E� �E� �E� �E� �E���E��E���E���E���E���E���E���E���E��E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E���E���E���E���E���E���E���E���E���E���E� �E� �E� �E� �E� �E� �E� �E׀�= � t�xP��!�E���E��E�M��M؋U�U��}��  4�}��  ��  �E����E��}��   ��  �M���8��$����E�-�  �E��}���  �M��$���E�   �E�h��U��]��E� �]��M��]ȍU�R�U؃���u�(���� "   �E�E���c  �E�   �E�h��M��]��U��]��E� �]ȍM�Q�U؃���u�ܨ��� !   �U�E���  �E�   �E�`��E� �]��M��]��U��]ȍE�P�U؃���u萨��� "   �M�E����  �E�   �E�`��U��]��E� �]��M��]ȍU�R�U؃���u�D���� !   �E�E���  �E�   �E�\��M��]��U��]��E� �]ȍM�Q�U؃���u������ "   �U�E���3  �E�   �E�\��E� �]��M��]��U��]ȍE�P�U؃��M�E����  �E�   �E�X��U�����  �E�   �E�X��E� �]��M��]��U��]ȍE�P�U؃���u�U���� "   �M�E���  �E�   �E�X��U��]��E� �]��M��]ȍU�R�U؃��E�E���S  �E�   �E�X��M��]��U��]��E� �]ȍM�Q�U؃���u�̦��� "   �U�E���  �E�   �E�X��E� �]��M��]��U��]ȍE�P�U؃���u耦��� !   �M�E���  �E�   �E�X��U��]��E� �]��M�����U��E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���O  �E�   �E�P��U��]��E� �]��M��]ȍU�R�U؃���u�ȥ��� !   �E�E���  �E�   �E�H��M��]��U��]��E� �]ȍM�Q�U؃���u�|���� !   �U�E���  �E�   �E�@��E� �]��M��]��U��]ȍE�P�U؃���u�0���� "   �M�E���k  �E�   �E�h��U�����E��M��]��U��]��E� �]ȍM�Q�U؃���u�Ԥ��� !   �U�E���  �E�   �E�`��E� ����M��U��]��E� �]��M��]ȍU�R�U؃���u�x���� !   �E�E���  �E�   �E�\��M�����U��E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���W  �E�   �E�8��U�����E��M��]��U��]��E� �]ȍM�Q�U؃���u������ !   �U�E����  �E�   �E�0��E� ����M��U��]��E� �]��M��]ȍU�R�U؃���u�d���� !   �E�E���  �E�   �E�(��M�����U��E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���C  �E�   �E�X��U��]��E� �]��M��]ȍU�R�U؃���u輢��� !   �E�E����  �E�   �E� ��M�����U��E� �]��M��]��U��]ȍE�P�U؃���u�`���� !   �M�E���  �E�   �E�H��U��]��E� �]��M��]ȍU�R�U؃���u����� !   �E�E���O  �E�   �E�P��M��]��U��]��E� �]ȍM�Q�U؃���u�ȡ��� !   �U�E���  �E�   �E���E� �M�M��U��]��E� �]��M��]ȍU�R�U؃���u�o���� !   �E�E���   �E�   �E���M��M�U��E� �]��M��]��U��]ȍE�P�U؃���u����� !   �M�E���T�E�   �E���U��M�E��M��]��U��]��E� �]ȍM�Q�U؃���u������ !   �U�E���M�3��@�����]�;���Ӟ�k����Z������/����3�� 	
�I ۢ7����K����O����@��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E���#`�l�l]������������������̋�U��j
�"�l3�]����������̋�U���h��  �(�P�)������E��M���  ���  ��   ���E�$�T������E�}� ~C�}�~�}�t�5h��  �U�R�ׅ�����E��   �E�P���E�$j������   �M�Q�E������$���E�$jj�Zz�����}���E�$�.�����]��E��E������Dzh��  �U�R�U������E��D�B�E��� th��  �M�Q�5������E��$�"�U�R���E��$���E�$jj��y������]������������������������������������������������������������������������������������̋�U��j
�"�`3�]����������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    j�j|�����E�    �E�x ��   �(��M��E�$���U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�(������/�M�M��U�z uh �j jXhp�j�<z������u�랋M�QR�������E�@    �E������   �j蠌����ËM�d�    Y_^[��]������������������������������������������������������������������������̋�U��j�h8�h)d�    P���SVW���1E�3�P�E�d�    �E�x �L  h (  h�9h	&j �M��	Qj �0������E�}� u3��   �U�R�h}�����E��E��M����M���v�U�U���� u�M�M�� ��j�z�����E�    �U�z ��   j�}�����E܃}� ��   �E���P�}�����E؋M�U؉Q�}� t[j h�   hp�h��h8��E�P�M���Q�U�BP蔙����P�C������M܋U�B��M܋U�B�A�M�U܉Q��E�P�������M�Q�$������E������   �j車����ËU�B�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������̋�U��j�hX�h)d�    P���SVW���1E�3�P�E�d�    j�
y�����E�    �E�x ��   �(��M��E�$���U��U�}� tY�E�M�;Qu�E��M�Q�P�E�P�������2�M�M��U�z u!h �j h�   hp�j��v������u�뛋M�QR谈�����E�@    �E������   �j�=�����ËM�d�    Y_^[��]���������������������������������������������������������������������̋�U���E��u	� (  f�M�URh�9h	&�EP�MQ�UR�������]���������������������̋�U��j�hx�h)d�    P���SVW���1E�3�P�E�d�    �E�x �a  j�]w�����E�    �M�y �*  h (  j �U��	Rj ��o�����E�}� u"�E�    j��E�Ph���6w�����E��  �M�Q�y�����E��U��E����E���v�M�M���� u�E�E��  ��j�Js�����E܃}� ��   �E�    �M���Q�'s�����E؃}� taj h4  hp�h��h(��U�R�E���P�M�Q�ؕ����P臃�����U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P�k������M�Q�_������E������   �j�������ËU�B�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    j�:u�����E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P�>������M�Q�2��������E������   �j�ǅ����ËM�d�    Y_^[��]������������������������������������������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y���������������������������������������������������������������������������������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������������������������������������������������������̋�U��j ��!]�����������������̋�U���"]� ����������������̋�U��EP�0�Q�"��]� �������������������̋�U��,�]����̋�U��Q�0�P�"�E��}� u �4�Q��!�E��U�R�0�P�"�E���]������������������������������̋�U��EP�MQ�8�R��!��]� ���������������̋�U���hd��"�E��}� u�|��3���  hX��E�P��!�0�hH��M�Q��!�4�h8��U�R��!�8�h,��E�P��!�<��=0� t�=4� t�=8� t	�=<� u,�0�6�"�4��"�8��"�<��"�0��=0��t�4�Q�0�R�"��u3���   �Nt���0�P��!�0��4�Q��!�4��8�R��!�8��<�P��!�<�������u��z��3��   h�7�0�Q��!�У,��=,��u	�z��3��rh  h��jh  j�Č�����E��}� t�U�R�,�P�8�Q��!�Ѕ�u	�gz��3��(j �U�R��������!�M���U��B�����   ��]������������������������������������������������������������������������������������������������������������������������������������̋�U��=,��t�,�P�<�Q��!���,������=0��t�0�R�"�0������1���]����������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    hd��"�E�E�@\� �M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@h �j��m�����E�    �M�QhR�"�E������   �j�~�����j�m�����E�   �E�M�Hl�U�zl u�E���Hl�U�BlP�������E������   �j�2~����ËM�d�    Y_^[��]��������������������������������������������������������������������������̋�U����$"�E��,�P�Hd���ЉE��}� u}j h�  h��jh  j�jm�����E��}� tW�M�Q�,�R�8�P��!�Ѕ�t%j �M�Q��������!�U���E��@�����j�M�Q��}�����E�    �U�R� "�E���]�����������������������������������������������������������̋�U��Q��d���E��}� u
j覄�����E���]�����������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P�}�����M܃y, tj�U܋B,P�}�����M܃y4 tj�U܋B4P��|�����M܃y< tj�U܋B<P��|�����M܃y@ tj�U܋B@P�|�����M܃yD tj�U܋BDP�|�����M܃yH tj�U܋BHP�|�����M܁y\� tj�U܋B\P�c|����j�j�����E�    �M܋Qh�U��}� t%�E�P�("��u�}� �tj�M�Q�|�����E������   �j�C{�����j�Ij�����E�   �U܋Bl�E�}� t4�M�Q�E������U�;�t�}� �t�E�8 u�M�Q��������E������   �j��z�����j�U�R�{�����M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��=,��tO�} u)�0�P�"��t�,�Q�0�R�"�ЉEj �,�P�8�Q��!�ЋUR�w���=0��tj �0�P�"]������������������������������������������̋�U����!]���̋�U���,"]���̋�U��Q�EP�MQ�UR���P�MQ�{�����E��E���]������������������̋�U��j j j�EP�MQ��z����]�������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�D   ���E��}� u�}� t�م����t
�Ѕ���M���E���]������������������������̋�U��Q�EP�MQ�UR�EP�MQ�   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP�Nw������u�} t	�M�   3��뗋�]�����������������������������̋�U��j j j�EP�s����]�������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�f�����E�    �=d� vU�d���9L�u6�p�����u!h�j h  h��j�d������u��L�    ��L����L��@��E؃=D��t�M�;D�u̃=P� tu�UR�EP�M�Q�UR�EPj j�P�����uP�} t%�MQ�URhP�j j j j �e������u�� h(�h��j j j j ��d������u��D  �U����  ��t�8���u�E�   �}�v3�MQh��j j j j�d������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h��h��j j j j�Dd������u̋M��$�MԋU�R�H������E܃}� u�} t	�E�    �r  �@����@��}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+D�;Mv�D�U�D��
�D������\�E�\��\�;P�v�\��P��=T� t�T��M܉H�	�U܉H��E܋T���U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉T�j�H�R�E܃�P��b����j�H�Q�U�E܍L Q�b�����UR�K�P�M܃� Q�b�����U܃� �U��E������   �j�/t����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�(������E��}� u�}� t������t
�����U���E���]����������������������������̋�U��Q�} v�����3��u;Es����    3��K�E�E�E�MQ�UR�EP�MQ���R�EP��������E��}� t�MQj �U�R�`�����E���]���������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�a�����E��}� u�}� t��~����t
��~���M���E���]������������������������̋�U��Qj j j�EP�MQ�UR�W�����E��E���]����������������������̋�U��j�h8�h)d�    P���SVW���1E�3�P�E�d�    j�:`�����E�    j�EP�MQ�UR�EP�MQ�b   ���E��E������   �j��p����ËE�M�d�    Y_^[��]����������������������������������������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�W�����  �} t�}� u�EP�MQ�q����3��  �=d� vV�d���9L�u6�3�����u!h�j h�  h��j�m]������u��L�    ��L����L��@��U�=D��t�E�;D�u̃=P� ty�MQ�UR�E�P�MQ�U�R�EPj�P�����uR�} t%�MQ�URh��j j j j ��]������u�� hx�h��j j j j �]������u�3��  �}��v`�} t)�UR�EP�M�Qh(�j j j j�o]���� ��u���E�Ph��j j j j�N]������u��|���    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh��j j j j��\������u�� h��h��j j j j��\������u��Qj�I�R�E�����P�  ����t1�MQhh�j j j j�\������u��X{���    3��t  �EP�^������u!h�j h  h��j�\[������u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!hh�j h#  h��j�[������u��d�M�Q����  ��u�E%��  ��u�E   �M�D�;Qs1�EPh(�j j j j�[������u��lz���    3��  �} t%�U���$R�E�P�]�����E��}� u3��_  �#�M���$Q�U�R��~�����E��}� u3��:  3�u��@����@��}� u|�=D��s9�U�D�+B�D����+D�;M�v�D�U��D��
�D������E��\�+H�\��\�U��\��\�;P�v�\��P��U��� �U�E��M�;Hv$�U��E�+BP�K�Q�U��E�BP�\Z����j�H�Q�U�U�R�CZ�����}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!h��j h�  h��j�Y������u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8�H�;M�t!ht�j h�  h��j�X������u̋E��H�H��U��z t�E��H�U����7�T�;M�t!h4�j h�  h��j�dX������u̋E���T��=T� t�T��E��B�	�M��H��U�T���M��A    �U��T��E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es�v���    3��g�E�E�E��} t�MQ�c�����E��UR�EP�MQ�U�R�EP�p�����E�}� t �M�;M�s�U�+U�Rj �E�E�P�V�����E��]����������������������������������������������������̋�U��Qj j j�EP�MQ�p�����E��E���]����������̋�U��j�hX�h)d�    P���SVW���1E�3�P�E�d�    3��} ���E��}� u!h�j h�  h��j�U������u̃}� u-��t���    j h�  h��h��h���l����3��c�}�v�t���    3��Nj�oV�����E�    j �UR�EP�MQ�UR�EP�������E��E������   �j�g����ËE�M�d�    Y_^[��]�������������������������������������������������������������������̋�U��j�EP�_����]�����������̋�U��j�hx�h)d�    P��SVW���1E�3�P�E�d�    j�zU�����E�    �EP�MQ�"_�����E������   �j�:f����ËM�d�    Y_^[��]����������������������������������̋�U��Q�=d� vU�d���9L�u6��v����u!h�j h  h��j�%S������u��L�    ��L����L��} u�l  �}uOj�I�P�M�����Q�	  ����t/�URh��j j j j�S������u��sr���    �  �=P� tDj j j �MQj �URj�P�����u%h��h��j j j j �RS������u���  �MQ��T������u!h�j h*  h��j�,R������u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!hX�j h0  h��j��Q������u̋8����m  j�H�P�M���Q�k  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ����Ph��j j j j�:R����(��u��<�U��� R�E��HQ�U��B%��  ����Qh��j j j j��Q���� ��u�j�H�P�M��Q�E��L Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ����Ph�j j j j�Q����(��u��<�U��� R�E��HQ�U��B%��  ����Qhx�j j j j�BQ���� ��u̋E��xue�M��y����u	�U��z t!h��j hi  h��j�P������u̋M��Q��$R�J�P�M�Q��P�����U�R��a�����Q  �E��xu�}u�E   �M��Q;Ut!h��j hw  h��j�O������u̋M��\�+Q�\��8�����   �M��9 t�U���M��Q�P�6�H�;E�t!hd�j h�  h��j�?O������u̋U��B�H��M��y t�U��B�M����5�T�;E�t!h0�j h�  h��j��N������u̋U���T��M��Q��$R�J�P�M�Q�O�����U�R�`�����(�E��@    �M��QR�J�P�M��� Q�iO������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�EP�S����]�����������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!h�j h�  h��j��L������u̃}� u1�|l���    j h�  h��h0�h��|d��������8  �=d� vV�d���9L�u6�p����u!h�j h�  h��j�NL������u��L�    ��L����L�j��M�����E�    �UR�N������u!h�j h�  h��j��K������u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!hX�j h�  h��j�K������u̋E��xu�}u�E   �M��Q�U��E������   �j��]����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������̋�U��Q�D��E��M�D��E���]������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    j�
L�����E�    �EP��L������te�M�� �M�U�B%��  ��tC�M�yt:�U�B%��  ��t*�M�yt!hX�j h?  h��j��I������u̋E�M�H�E������   �j�e\����ËM�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�P��E��M�P��E���]������������������̋�U��P�]����̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�����������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �8���u
�   ��  j�FJ�����E�    �K���E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$�8�h��h��j j j j �(I������u��   h��h��j j j j �I������u��dh��h��j j j j ��H������u��Bhx�h��j j j j �H������u�� hD�h��j j j j �H������u��E�    ��  �E�   �T��E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  �����U���E�8�j�H�P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh��j j j j �G����(��u��-�E�� P�M�QR�E�Ph��j j j j �G���� ��u��E�    j�H�R�E�H�U�D
 P�2�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph�j j j j �G����(��u��-�U�� R�E�HQ�U�Rhx�j j j j ��F���� ��u��E�    �M�y ��   �U�BP�J�Q�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� Rhx�j j j j �wF���� ��u��"�M�� Qh��j j j j �SF������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rh��j j j j �F����(��u��-�M�QR�E�� P�M�QhL�j j j j ��E���� ��u��E�    �G����E������   �j�VW����ËE܋M�d�    Y_^[��]ÍI �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �8��E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!hH�j hy  h��j��B������u̃}� u0�b���    j hy  h��h �hH��Z�����8��sj�[D�����E�    �8��M�}�t7�U��t�d�   ��E��%��  �d��L�    �M�8��E������   �j��T����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    3��} ���E��}� u!hT�j h�  h��j�yA������u̃}� u+�,a���    j h�  h��h�hT��,Y�����s�8���u�fj��B�����E�    �T��E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j�mS����ËM�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��3��} ��]����������������̋�U��} u3��1j j �E�� P��I������u3���M�� Qj ���R�0"]������������������������������̋�U��j�h8�h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP�B������u3���   j�A�����E�    �M�� �M��U��B%��  ��t"�M��yt�U��B%��  ��t	�M��yukj�UR�EP��H������tU�M��Q;UuJ�E��H;@�<�} t�U�E��H�
�} t�U�E��H�
�} t�U�E��H�
�E�   ��E�    �E������   �j�+Q����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U��Q�EP�@������u�����M�� �M��U��B��]������������������̋�U��Q�X��E��M�X��E���]������������������̋�U��X�]����̋�U��j�hX�h)d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!h�j h�  h��j�9=������u̃}� u.��\���    j h�  h��h��h���T�����m  j�>�����E�    �U�T���E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡT��E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�Rh��j j j j ��<���� ��u���M�Qhp�j j j j �<������u������E�P��H,�U�D��B0�E������   �j�0N����ËM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E�}� u!h�j h�  h��j�:������u̃}� u0�nZ���    j h�  h��h��h��nR����3��  3҃} �U��}� u!h\�j h�  h��j�R:������u̃}� u0�Z���    j h�  h��h��h\��R����3��0  3Ƀ} ���M�}� u!h4�j h�  h��j��9������u̃}� u0�Y���    j h�  h��h��h4��Q����3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u�8���t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M���E���M��7��P�MQ�#   ���M��X����]��������������������̋�U��j�hx�h)d�    P���SVW���1E�3�P�E�d�    �E�    j�s9�����E�    h��h��j j j j �8������u̃} t�M��U�T��E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�8���u��  �U�z twj j�E�HQ��@������tj�U�BP�4"��t$�M�QRh��j j j j ��7������u��)�M�QR�E�HQh��j j j j �7������u̋E�HQhx�j j j j �}7������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph8�j j j j �/7���� ��u̃=X� t,j�U�� R�4"��u�E�HQ�U�� R�X�����E�P�MQ�  ���   �U�zu;�E�HQ�U�� Rh�j j j j �6������u̋M�Q�UR�x  ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Ph��j j j j �W6���� ��u̋U�R�EP�  ��������E������   �j��G�����h��h��j j j j �	6������u̋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���t���3ŉE��EP�M���A���E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M��3����t3�M��3������   ~ �M���2��PhW  �E�P�hM�����E��hW  �M�Q�M���2��P�E-�����E��}� t	�U��U���E�    �E��M��L��S����U��S���     �E�Ph���M�k��1   +�R�E�k��L�Q�F������}*j h	  h��h��h��j"j�R���R��-���� �R���M��������U��D� �E�P�M�Qh��j j j j �3������u̍M��CS���M�3���U����]������������������������������������������������������������������������������������������������������������������̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP�RI���E]������������������̋�U���8���3ŉE��E�P�h8�����}� u�}� u�8���t7�}� t1h �h��j j j j �s2������u�j �J�����   �3��M�3��T����]������������������������������������̋�U���3��} ���E��}� u!h�j h�	  h��j�1������u̃}� u.�P���    j h�	  h��h��h��H�����   �E�    �	�U����U��}�}>�E�����Q�U��E�L�Q�U��E�L�Qh��j j j j �k1���� ��u�볋E�H,Qhd�j j j j �G1������u̋E�H0Qh<�j j j j �%1������u̋�]�������������������������������������������������������������������̋�U��j j j �EP�MQ�?1����]�������������������̋�U��EP�MQj �UR�EP�1����]���������������̋�U��j j j �EP�MQ�UR�T0����]���������������̋�U��j j j �EP�MQ�UR�EP�:����]�����������̋�U��EP�MQj �UR�EP�MQ��/����]�����������̋�U��EP�MQj �UR�EP�MQ�UR�4:����]�����������������������̋�U��j j �EP�MQ�UR�0����]�����������������̋�U���(�E��#E������E�u!hl�j h�
  h��j�P.������u̃}� u0�N���    j h�
  h��h,�hl��F����3��@  �} t�U;Ur	�E�    ��E�   �E܉E��}� u!h��j h�
  h��j��-������u̃}� u0�M���    j h�
  h��h,�h���E����3��   �}v�U�U���E�   �E؃��E3�+M���M�U�E�L�M��UU��U�E;E�v�M���    3��i�MQ�URj�E�P� '�����E�}� u3��F�M�M�M�U��#�+M�M��E�+E���E�j�I�Q�U���R�-�����E��M��E���]������������������������������������������������������������������������������������������������������������������������̋�U��j j �EP�MQ�UR�EP�"-����]�������������̋�U��j j �EP�MQ�UR�EP�MQ�f7����]���������̋�U���4�} u!�EP�MQ�UR�EP�MQ�@-�����  �} u�UR�AL����3��  �E������E�j�H�Q�U��R�V�������t1�EPh(�j j j j�^,������u��'K���    3��C  j�I�R�E���P��������u�MQh��j j j j�,������u̋E��#E������E�u!hl�j h�  h��j��*������u̃}� u0�J���    j h�  h��h��hl��B����3��  �} t�U;Ur	�E�    ��E�   �EԉE؃}� u!h��j h�  h��j�i*������u̃}� u0�J���    j h�  h��h��h���B����3��  �U��P�7�����M��U++E�}v�E�E���E�   �MЃ��M3�+U���U�E�M�T�U�EE�E�M;M�v�I���    3��   �UR�EPj�M�Q�|#�����E��}� u3��   �U�U�U�E��#�+U�U��M�+M���M�j�I�R�E���P�4*�����M��U���E�;Ev�M�M���U�ŰE�P�MQ�U�R�A6����j�E��Q�v<�����E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es��G���    3��s�E�E�E��} t�MQ�UR�EP�A�����E��M Q�UR�EP�MQ�U�R�EP�(�����E�}� t �M�;M�s�U�+U�Rj �E�E�P�s(�����E��]��������������������������������������������������������̋�U��EP��G����]�������������̋�U��Q�} u�   �E������E�j�H�Q�U��R���������t!�EPh��j j j j��'������u��Lj�I�R�E���P��������u�MQh��j j j j�'������u�j�E��Q��9������]�����������������������������������������������������̋�U��Q�<��E��M�<��E���]������������������̋�U��Q�`��E��E���]�����������̋�U��`�]����̋�U��EP�MQ�UR�}#����]���������������������̋�U��� �E�    �E�    �E�    �E�    �E�    3��} ���E�}� u!h�j h�  h��j�p%������u̃}� u.�#E���    j h�  h��h��h��#=��������w�E�    �U������U��E��Q�2�����E��U��E+�E�3�+M���M�}v�U�U���E�   �E����E�M�U�D
+E�E�M�+M�+M�M��E���]�������������������������������������������������������������������̋�U��Q�=�� th���>������t�EP�������5��h4�h��sD�����E��}� t�E��Gh�#�n$����h�h ��R  ���=\ th\�'>������tj jj �\3���]���������������������������������������������������̋�U��j j �EP�>  ��]���������̋�U��j j�EP�  ��]���������̋�U��jj j �   ��]�����������̋�U��jjj ��  ��]�����������̋�U���<���EP�'����h�   �&��]��������������̋�U��Q����E��	�M����M��}� t�U��: tj�E��Q�!6������j���R�6�������    ����E��	�M����M��}� t�U��: tj�E��Q��5������j���R��5�������    j�|�P�5����j�x�Q�5����j�TR��!P�}5�����|�    �x�    �:*���T�H�P�("��u'�=H� �tj�H�Q�25�����H� ��H�R�"��]�����������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �^6���E�    �=���U  ���   �E����} ��   �TQ��!�E�}� ��   �PR��!�E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�(���U�9u��E�;E�s�h�M؋R��!�E��(���M؉�U܋TR��!�EСPP��!�E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���hL�h8��A  ��hT�hP��/  ���=�� u#j��1������ t���   �B���v1���E������   ��} t��B��Ã} t����   ��B���MQ�m#�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������̋�U���h@��"�E��}� th,��E�P��!�E��}� t�MQ�U���]�����������������̋�U��EP�B�����MQ�8"]�������������������̋�U��j� ����]���������������̋�U��j��0����]���������������̋�U��Q�S&���E��E�P��?�����M�Q��:�����U�R�*�����E�P�������M�Q�l!�����U�R�*������]����������������������̋�U��E;Es�M�9 t�U��ЋM���M��]�����������������������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�����������������̋�U���3��} ���E��}� u!h �j h�  h��j��������u̃}� u0�<���    j h�  h��h��h ��4�����   �y3҃=�� �U��}� u!h\�j h�  h��j�������u̃}� u0�:<���    j h�  h��h��h\��:4�����   ��M����3���]������������������������������������������������������������������̋�U���3��} ���E��}� u!h �j h�  h��j��������u̃}� u0�v;���    j h�  h��hl�h ��v3�����   �y3҃=�� �U��}� u!hD�j h�  h��j�W������u̃}� u0�
;���    j h�  h��hl�hD��
3�����   ��M����3���]������������������������������������������������������������������̋�U���p�E�P�L"h�   h��jj@j �k9�����E��}� u�����  �M��@��    �	�U���@�U��@   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M���;U���   h�   h��jj@j �H8�����E��}� u���E��   �M��U���@���� ���	�M���@�M��U���@   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R�H"��t[�E����M������@�M��U��E���
�U��E���Jh�  �U���R�D"��u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M���@�M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P�@"�E��}����   �}� ��   �M�Q�H"�E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�D"��u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A�������R�<"3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �	�E����E��}�@}y�M��<�@ tg�U���@�E��	�M���@�M��U���@   9E�s�M��y t�U���R�P"��j�E���@Q�(�����U���@    �x�����]���������������������������������������������������̋�U����=X u�8���E�    ����E��}� u����e  �M����t,�E����=t	�U����U��E�P������M��T�U���juh��jj�E���P�"3�����E�M����=�� u�����   ����U��	�E�E��E��M������   �E�P�G�������E��M����=��   j~h��jj�E�P�2�����M��U�: uj���P�!'�������    ����rj h�   h �h�h���M�Q�U�R�E�Q�4����P�P"�����U���U��B���j���P�&�������    �M��    �@   3���]��������������������������������������������������������������������������������������������������������������������̋�U����E�    �=X u�p6����� h  h��j �T"h����6�����=� t�����t���U���E���E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   h��j�M��U���P�������E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�   ���U����t��E��x�3���]�������������������������������������������������������������������������̋�U��E���]�����������������̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�#������t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P�$!������t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R�� ������t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �\"�E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j ��!�E��}� tjJh j�M�Q�H�����E�}� u�U�R�X"3��Dj j �E�P�M�Q�U�R�E�Pj j ��!��uj�M�Q������E�    �U�R�X"�E��]������������������������������������������������������������������������̋�V�����=��s���t�Ѓ�����r�^����������̋�V� ���=p�s���t�Ѓ���p�r�^����������̋�U��Q�E�   j h   j �`"����=�� u3���   ��]�������������������������̋�U����P�d"���    ]�������������������̋�U��=�� uh� j jhhH j��
������u̡��]�������������̋�U���0�E� �E�   �E���E��M����M�U��B3���EԋM�Q�U�R��  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M�����E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=�� t h����#������tj�UR������M����U��$���E��H;M�th���U�R�M����U��S���E��M�H�U�R�E�P��   ���U�M�I��+�������&�U��z�th���E�P�M������������E��M߅�t�U�R�E�P�   ���E��]������������������������������������������������������������������������������������������������������������������������̋�U����E�8�t%�M��E��M��U�EB3E��E��M��+���M�Q�E��M��U�EB3E��E��M��y+����]���������������������������������̋�U����E�    �E�    �=��N�@�t���%  ��t����щ���   �U�R�t"�E��E�M�3M��M��p"3E�E���!3E�E��l"3E�E�U�R�h"�E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M����U��҉����]����������������������������������������������������������������̋�U��}csm�u�EP�MQ�!������3�]����������̋�U����\���E��}� u3���  �E��H\Q�UR�S  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  �h�U��	�E����E��hl9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��;Ut�E����E��tk�M9M�s�ڋtk�U9U�s
�E��;Mt3���E���]������������������������̋�U���(  � �����������5���=��f��f��f���f���f�%��f�-������E ���E���E���������P�  �������	 ����   ��������������������!�H�j�����j ��"h���"�=H� u
j�����h	 ��|"P�x"��]����������������������������������������������������������������������������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh�j jphj�������u̃}� u.�!���    j jphh�h����������)  �} t�} u	�E�    ��E�   �M̉MЃ}� uh�j jshj�������u̃}� u.�;!���    j jshh�h��>��������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�i�����E��} u�E��P�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �������EċE���]�������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�$����]���������������̋�U��=�� u0�EP���E�$�����$���E�$�MQj�i����$�!��y��� !   h��  �UR�:	�����E]���������������������������������̋�U����E�E�]��=�� u1�EP���E��$���E�$���E�$�MQj������$�!������ !   h��  �UR������E���]����������������������������������̋�S�܃������U�k�l$���   ���3ŉE��C P�KQ�SR�������u)�E�����E��KQ�SR�CP�KQ�S R�E�P�%�����KQ��������|����=�� u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q������$�%���|���R�����h��  �C P������C�M�3��U!����]��[��������������������������������������������������������������������������̋�S�܃������U�k�l$���   ���3ŉE��C(P�K Q�SR��������u;�E����E��M������M��C�]��S R�CP�KQ�SR�C(P�M�Q�������SR�������|����=�� u?��|��� t6�C(P���C �$���C�$���C�$�KQ��|���R�����$�%���|���P�����h��  �K(Q�O�����C �M�3�� ����]��[�����������������������������������������������������������������������̋�U����E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U�������������M�Q���ЋE�P�M�����҃������E�H���ʋU�J�E�����Ƀ������U�B�����M�A�U�������������M�Q���ЋE�P�M��� ��҃����E�H���ʋU�J����E��E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E���t�M�Q���E�P�M��� t�U�B���M�A�U�%   �E�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�M����E��1�M�������E���M�������E���M�����E��M���   �U�t5�}�   t�}�   t�1�E����U�
�"�E������U�
��E������U�
�E%�  ���M��� ��ЋE��}  tT�M�Q ���E�P �M�Q ���E�P �M�U��Y�E�H`���U�J`�E�H`���U�J`�E�M��XP�X�U�B ���M�A �U�B �����M�A �U�E� �Z�M�Q`���E�P`�M�Q`�����E�P`�M�U��YP����EPjj �M�Q��!�U�B����t�M�����E��M�Q����t�E�����U�
�E�H����t�U�����M��U�B���t�M����E��M�Q��t�E���ߋU�
�E����M�}�wb�U��$��0�E���������   �U�
�@�E���������   �U�
�(�E���������   �U�
��E��������U�
�E������M�t�}�t�}�t.�;�U�%����   �M��%�U�%����   �M���U�%�����M��}  t�U�E�@P���M�U�BP���]�0�/�/�/�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR� ����]�����������������������̋�U��j�EP�MQ�UR�EP�MQ�UR�R ����]�����������������������̋�U���D�E���E��M��t �U��tj�f�����E�����E��  �M��t �U��tj�>�����E�����E��s  �M���   �U���  j������E%   �E��}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z����]��������]؋U�E���   �E�������z����]��������]ЋM�E���Z�U�������z����]��������]ȋE�E���,�M�������z����]��������]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�E������]�M��   �M��}�����}�E��H��]��E�   �   ���]�����Au	�E�   ��E�    �U��U��E��f�E��M��f�M��	�U����U��}����}:�E��t�}� u�E�   �M���M�U��t�E�   ��E�M���M�봃}� t�E����]�U�E����E�   �}� t
j�������E�����E��M��t�U�� tj ������E����E�3��}� ����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �EP�  ���E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R��������E�P�������u�MQ�������E��"� h��  �U(R�������EP��������E ��]�������������������������������������������������̋�U��Q�E�E��}�t�}�~ �}�~��W��� !   ��J��� "   ��]��������������������̋�U��Q�E�    �	�E����E��}�}�M��͠�;Uu�E��Ť����3���]�������������������������������̋�U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]���������������������������������������̋�U����E�]��E�  �E��M���  �U����f�M��E���]��������������������������̋�U��Q�E%�  ��f�E��M����  f�M��E���]��������������������̋�U���E%�  ���ȋU�����P���E�$�����]��������������̋�U����E�]��E%�  �M���f�E��E���]����������������������̋�U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]�������������������������������������������̋�U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U�U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$������]��.j ���E�$������]��U���  ����-�  �E��M�U���E���]�������������������������������������������������������������������������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]������������������̋�U����E��t
�-���]���M��t����-���]������U��t
�-���]���E��t	�������؛�M�� t���]����]�������������������������̋�U��Q�=` t�]���E�    �E���]�������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �e�=` ��   �E��@tp�= � tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe�� �    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]�������������������������������������������������������̋�U��Q�=` t�]��e���U���]�����������������̋�U��Q�=` t� ����E��E���?�E���E�    �E���]����������������̋�U��Q�=` t������E��E���?�E�������E�    �E���]���������������������������̋�U����=` t8�����E��E#E�M��#M���E��U������U��U��E�P��������E�    �E���]�������������������������̋�U��Q�)����E��E��?E��E��M�Q�2�������]�����������������������U���0���S�ٽ\�����=�� t�V�����8����   [����ݕz������U���U���0���S�ٽ\����=�� t������8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���������   [�À�8�����=�� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �X�����������H����s4�h�,ǅr���   �P�����������@����v�`VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P������_^�E�����U���0���S�u�u�   ���ٽ\�����8�����7�������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[������������������������������������������������������������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp��������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-���p��� ƅp���
��
�t������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    ����t
j
�-������s����E��}� t
j����������tjh  @j�d�����j������]��������������������������������̋�U��Q���E��M��#M��U#Uʉ��E���]���������������������̋�U��j���������tj���������u#�=�uh�   �V�����h�   �I�����]�������������������������̋�U��Q�E�    �	�E����E��}�s�M��U;��u�E�������3���]�������������������������������̋�U���   ���3ŉE�EP�]������E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j�g����������������� t������t���E�   ��E�   �}� ��  j��������tj����������   �=���   j��@"�E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P�������P������Q�U�R��"��  �}�   ��  ǅ������������-�����  +ȉ�����������������j h  h�h�h�h�h  h���� ����P�������3�������f��  h  ������Rj ��"��u:j h  h�h�hh�������P������Q� ����P�|�����������R�d���������<vk������P�M������������TA�������j h  h�h�hHjh<������+�������������+�Q������R�������P�������j h  h�h�h�h�h  h���a�����P�������j h  h�h�h��E�Ph  h���,�����P������h  h�h��������M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   ���3ŉE�}��  �E�E���p����M�ǅd���    ǅh����   ��h���R�E�P�MQ�UR�EP��������l�����l��� ��   �$"��zt�  j j �MQ�UR�EP�x�������h�����h��� u��   j^hxjj��h���Q��������E��}� u��   ǅd���   ��h���R�E�P�MQ�UR�EP��������l�����l��� u�   jihxjj��l���Q�f������U���E��8 u�]j jlh h�hP��l�����Q�U�R��l���P�M��R�>�����P��������d��� tj�E�P������3��-  ��d��� tj�M�Q�v���������  �  �}��   �U��\�����\����     j j �MQ�UR��"��`�����`��� u�Zh�   hxjj��`���P�w�������\������\����: u�(��`���P��\����R�EP�MQ��"��u�3��mj��\����P��������\����    ����I�D�} u>ǅX���    j��X���R�E    P�MQ��"��u�����U��X����3������M�3��R�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�$�]�����������������̋�U��E�U��DV�u�     j�E�P3�NVf�
��"��u3�^��]ËM�U�E�QRP��"��t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=,� u �=(� uH�  �(���t:�,���(�h�P��!3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�Rh�V�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ��"P��"�����   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ��"P��"�M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE��=-� t3��M�3��������]��-���   ����   VWh��"�= "�5�"��t?h  ������QP�օ�t,h  ������R������P��  ����t������Q�ׅ�uBh  ������Rj �օ�t,h  ������P������Q�  ����t������R�ׅ�u3�_^�M�3�������]����������������������������������������������������������������̋�U���  ���3ŉE�Vh�� "����u^�M�3�������]�W�=�!h�V�׉�������u_^�M�3��y�����]�Sh�V�׋؅�t4h�V�׋���t&������Pjj hHh  ���������tV��"[_3�^�M�3��#�����]Í�����Q������������R������Pj hQǅ����  �Ӌ�����R����V��"��u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M���������E��������H���P���H���Pf���Hf�P������P� "�M�[_3�^������]����������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE��EV�uh   ������Qh   ������Rh   ������Qj�U�RP�������$��t3�^�M�3��D�����]�h������j	P��������u�h������jQ��������u�������R������P�E������Q�U�RPV�����M������3�@^�������]��������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh�j jahxj���������u̃}� u.�y����    j jahxhDh��|���������h  3҃} �U؃}� uhj jbhxj�b�������u̃}� u.�����    j jbhxhDh����������  j��������E�    ���M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H��j�U�R��������43�uh�j jhxj�W�������u��E������	����    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;�tM�U�z t�E�H�U���M��E�H�J�U��    �E���H���E��M���h�   hljj�������E�}� u�E������X����    �L�U��    �E���H�=� t���E��M��A   �E�   �U�E�B�M���E������   �j�������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR�.�����]���������̋�U��P  �I������3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �T"��u8j h<  hxhlh�h�h  ������Q�^�����P�������������U��E�P�b�������@v]�M�Q�Q������U��D��E�j hE  hxhlh�j��Q�U�������+й  +�Q�U�R������P�������} t'�EP���������@v�MQ��������U�DÉE��U�����������H����     �}uǅ����8�
ǅ����+��U���t�M�������
ǅ����+��U���t�}uǅ����(�
ǅ����+��M���tǅ����$�
ǅ����+��} t�E�������
ǅ����+��} tǅ�����
ǅ����+��} t�M�������
ǅ����+��} tǅ�����
ǅ����+��}� t�U��������'�} t�E�������
ǅ����+��������������}� tǅ����0�
ǅ����+��} tǅ���� �
ǅ����+�������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U��\Ph�h�  h   ������Q�8�����D�E�}� }*j h`  hxhlh��j"j�A����R������ �1�����������}� }8j he  hxhlh�h�h   ������R�K�����P�������h  h�������P�@�����������������uj������j����������u�   �3��M�3��.�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh�j jahxj�V�������u̃}� u.�	����    j jahxh�h�����������h  3҃} �U؃}� uhj jbhxj���������u̃}� u.�����    j jbhxh�h����������  j�\������E�    ���M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H��j�U�R�e������43�uh�j jhxj���������u��E����������    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;�tM�U�z t�E�H�U���M��E�H�J�U��    �E���H���E��M���h�   hljj�������E�}� u�E�����������    �L�U��    �E���H�=� t���E��M��A   �E�   �U�E�B�M���E������   �j�U�����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP��������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR������]���������̋�U��X"  ��������3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj ��"��u8j h<  hxhd!h� h�h  ������R������P�������������E��M�Q�}�������@v`�U�R�l������M��TA��U�j hE  hxhd!h�j��P�M�������+����  +���P�M�Q������P�!������} t'�UR��������@v�EP��������M�TA��U������� ������������     �}uǅ������
ǅ������M���t�E�������
ǅ������M���t�}uǅ������
ǅ������E���tǅ������
ǅ������} t�U�������
ǅ������} tǅ������
ǅ������} t�E�������
ǅ������} tǅ������
ǅ������}� t�M��������'�} t�U�������
ǅ������������������}� tǅ����<�
ǅ������} tǅ����l�
ǅ�����������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M���Rh�h�  h   ������P觽����D�E�}� }*j h`  hxhd!h��j"j������Q������ ������������}� }8j hc  hxhd!h�h�h   ������P������P������h  h(������Q�z�����������������uj������j����������u�   �3��M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�D������E��E�    �E���]�����������������̋�U����E%�����E�M#M��������   �} tj j �J������U�3�t	�E�   ��E�    �M��M��}� uhH"j j1h�!j蔾������u̃}� u-�G����    j j1h�!h�!hH"�J������   �/�} t�EP�MQ辽�����U���EP�MQ觽����3���]����������������������������������������������������������������̋�U��E�0�]�����������������̋�U��Q�0��E��M�Q��!�E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�������]����������������������̋�U��jh �j������h ��|"P�x"]����������������������̋�U���8  ���3ŉE��}�t�EP������ǅ����    jLj ������Q谽�����������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M��������!�E�j ��"�U�R��"���������� u�}� u�}�t�EP�������M�3��)�����]�������������������������������������������������������������������������������������������������̋�U��Q�E�    �0��E��M�Q��!�E��UR��!�E�E�0��E���]������������������̋�U��Q�E�    �0��E��M�Q��!�E��E���]�����������������������̋�U��EP�MQ�UR�EP�MQ������]�������������̋�U��EP�MQ�UR�EP�MQ�����]����������������̋�U����EP�M��!����M�誹����t2�M�螹������   ~�M�苹��Ph  �UR��������E��h  �EP�M��c���P�ֳ�����E�M�M�M������E��]��������������������������������������������̋�U��=L� uh  �EP�v�������j �MQ������]�������������̋�U����EP�M��1����M�躸����t/�M�许������   ~�M�蛸��Pj�UR�������E��j�EP�M��y���P�������E�M�M�M������E��]����������������������������������̋�U��=L� uj�EP虴������j �MQ�]�����]����������������̋�U����EP�M��Q����M��ڷ����t/�M��η������   ~�M�軷��Pj�UR�+������E��j�EP�M�虷��P�������E�M�M�M�������E��]����������������������������������̋�U��=L� uj�EP蹳������j �MQ�n�����]����������������̋�U����EP�M��q����M��������t/�M���������   ~�M��۶��Pj�UR�K������E��j�EP�M�蹶��P�,������E�M�M�M�������E��]����������������������������������̋�U��=L� uj�EP�ٲ������j �MQ������]����������������̋�U����EP�M������M�������t2�M���������   ~�M������Ph�   �UR�h������E��h�   �EP�M��ӵ��P�F������E�M�M�M������E��]��������������������������������������������̋�U��=L� uh�   �EP��������j �MQ������]�������������̋�U����EP�M������M��*�����t/�M���������   ~�M�����Pj�UR�{������E��j�EP�M�����P�\������E�M�M�M������E��]����������������������������������̋�U��=L� uj�EP�	�������j �MQ������]����������������̋�U����EP�M�������M��J�����t/�M��>�������   ~�M��+���Pj�UR�������E��j�EP�M��	���P�|������E�M�M�M��<����E��]����������������������������������̋�U��=L� uj�EP�)�������j �MQ�n�����]����������������̋�U����EP�M�������M��j�����t2�M��^�������   ~�M��K���Ph  �UR�������E��h  �EP�M��#���P薭�����E�M�M�M��V����E��]��������������������������������������������̋�U��=L� uh  �EP�6�������j �MQ������]�������������̋�U����EP�M�������M��z�����t2�M��n�������   ~�M��[���PhW  �UR��������E��hW  �EP�M��3���P覬�����E�M�M�M��f����E��]��������������������������������������������̋�U��=L� uhW  �EP�F�������j �MQ�|�����]�������������̋�U����EP�M������M�花����t2�M��~�������   ~�M��k���Ph  �UR��������E��h  �EP�M��C���P趫�����E�M�M�M��v����E��]��������������������������������������������̋�U��=L� uh  �EP�V�������j �MQ������]�������������̋�U����EP�M������M�蚰����t/�M�莰������   ~�M��{���Pj �UR��������E��j �EP�M��Y���P�̪�����E�M�M�M������E��]����������������������������������̋�U��=L� uj �EP�y�������j �MQ������]����������������̋�U��}�   ���]��������������̋�U��E��]���̋�U��Q�EP�MQ��������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP��������u�}_t	�E�    ��E�   �E���]�������������̋�U��Q�EP�MQ�z�������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP���������u�M��_t	�E�    ��E�   �E���]�������������������������̋�U��E�� ]���̋�U���4�EP�M�������}   ��   �M��=�����t/�M��1�������   ~�M�����Pj�UR�������E��j�EP�M������P�o������Ẽ}� t,�M���������   �E��M��M������E��*  ��U�U܍M�������E��  �M�蠭��� ���   ~D�M�荭��P�M�����   Q��������t"�U�����   �U��E�E��E� �E�   ������� *   �M�M��E� �E�   j�M��+�����BPj�M�Q�U�R�E�Ph   �M��
�����QR�M������P�Կ����$�E�}� u�E�E؍M��)����E��A�}�u�M��MԍM������E��'��U��E���ЉUЍM�������E���M��������]����������������������������������������������������������������������������������������������������������������������������̋�U��Q�=L� u$�}A|�}Z�E�� �E���M�M��E���j �UR��������]���������������������������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    誷���E��E��Hp#H�t�U��zl ��   j跭�����E�    �E��Hh�M�U�;H�tI�}� t%�E�P�("��u�}� �tj�M�Q�#������U�H��Bh�H��M�U�R�"�E������   �j�*�������	�E��Hh�M�}� u
j ��������E�M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h8�h)d�    P���SVW���1E�3�P�E�d�    �E������S����E��0����E܋Hh�M��UR��  ���E�E��M;H�  hN  h�"jh   �k������E��}� ��  �U܋rh��   �}��E��     �M�Q�UR贬�����E؃}� ��  �E܋HhQ�("��u�U܁zh �tj�E܋HhQ聽�����U܋E��Bh�M܋QhR�"�E܋Hp���-  �H����  j葫�����E�    �E��H�D��U��B�H��M��Q�L��E�    �	�E���E�}�}�M�U�E�f�TPf�M8����E�    �	�E���E�}�  }�M�M�U�A��@����E�    �	�M���M�}�   }�U�U�E䊊  ��H��׋H�R�("��u�=H� �tj�H�P�[������M��H��U�R�"�E������   �j�m�������(�}��u"�}� �tj�E�P�������o����    ��E�    �E؋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��d�    P��$���3�P�E�d�    �E�    �E�P�M��[����E�    �4�    �}�u)�4�   ��"�E��E������M�� ����E��}�c�}�u)�4�   ��"�E��E������M�������E��N�4�}�u.�4�   �M��e�����Q�U��E������M������E���E�E��E������M������EЋM�d�    Y��]����������������������������������������������������������������������������̋�U���,���3ŉE�V�EP�������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0��P�;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E����`��M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E���L��UU��B��MM��A����v����U�E�B�M�A   �U�BP��  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��pT�f�DJ�ӋMQ�C  ��3��  �����} t!�}��  t�}��  t�UR��"��u����k  �E�P�MQ��"���9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�\  ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=4� t�EP�  ��3�����^�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���  �M��}�w-�U���؅�$�ą�  ��  ��  �	�  �3���]ÍI ���������� ������������������������������������̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U���<��A���E�    �	�M����M��}�   }�UU��E���=���  �׋�]���������������������������������������������������������̋�U���(  ���3ŉE�������P�M�QR��"���-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj 蛰���� j �M�QRh   ������Ph   ������Qh   �U�BPj 蟱����$j �M�QRh   ������Ph   ������Qh   �U�BPj �h�����$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3��������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��J����M��ӛ���H�y t �M�����P�B�E�M�������E����E�    �M������E���M��ۼ����]������������������������������������̋�U��=X uj��������X   3�]����������̋�U��Q�EP�"�M���    t�U���   P�"�M���    t�U���   P�"�M���    t�U���   P�"�M���    t�U���   P�"�E�    �	�M����M��}�m�U����E�|HL�t$�M����U�|
P t�E����M�TPR�"�E����M�|L t$�U����E�|T t�M����U�D
TP�"넋M���   �´   R�"��]���������������������������������������������������������������������������������̋�U��Q�} �  �EP�("�M���    t�U���   P�("�M���    t�U���   P�("�M���    t�U���   P�("�M���    t�U���   P�("�E�    �	�M����M��}�m�U����E�|HL�t$�M����U�|
P t�E����M�TPR�("�E����M�|L t$�U����E�|T t�M����U�D
TP�("넋M���   �´   R�("�E��]������������������������������������������������������������������������������������̋�U��Q�E���    ��   �M���   ����   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�߫�����M���   R英�����E���    t4�M���   �: u&j�E���   Q蟫�����U���   P������j�M���   R�y�����j�E���   Q�e������U���    to�E���   �9 uaj�U���   -�   P�2�����j�M���   ��   R������j�E���   ��   Q�������j�U���   P�������M���   P�t8�U���   ���    u&�M���   R�ʵ����j�E���   Q裪�����E�    �	�U����U��}���   �E����M�|HL�t:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP�:������M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h@#j h�   h�"j��������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ菩���������j�UR�|�������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�������}� t�E�P�د�����}� t�M��9 u�}� �t�U�R荹�����E��]������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    ������E��E��Hp#H�t	�U��zl uDj�������E�    ��P�M���lQ蓰�����E��E������   �j�æ������藟���Pl�U�}� u
j 脮�����E�M�d�    Y_^[��]�����������������������������������������������������������̋�U���@���3ŉE��E�    �E�    �EP�M��I����M��Ғ��Pj j j j �MQ�U�R�E�P�ת���� �E��MQ�U�R蒴�����E��E���u8�}�u�E�   �M��ϳ���E��j��}�u�E�   �M�賳���E��N�:�M���t�E�   �M�蕳���E��0��U���t�E�   �M��w����E���E�    �M��c����E��M�3�������]�������������������������������������������������������������������������������̋�U��j �EP�MQ�u�����]�������̋�U���@���3ŉE��E�    �E�    �EP�M��ٟ���M��b���Pj j j j�MQ�U�R�E�P�g����� �E��MQ�U�R�c������E��E���u8�}�u�E�   �M��_����E��j��}�u�E�   �M��C����E��N�:�M���t�E�   �M��%����E��0��U���t�E�   �M������E���E�    �M������E��M�3�觴����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�������]�������̋�U���@���3ŉE��E�    �E�    �EP�M��i����M�����Pj j j j �MQ�U�R�E�P������� �E��MQ�U�R�ڱ�����E��E���u8�}�u�E�   �M������E��j��}�u�E�   �M��Ӱ���E��N�:�M���t�E�   �M�走���E��0��U���t�E�   �M�藰���E���E�    �M�胰���E��M�3��7�����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�E�����]�������̋�U����E�E��M�Q�U�3��} ���E�}� uh,�j j7h�)j�'�������u̃}� u0�ڮ���    j j7h�)h�)h,��ݦ�����   �$  3�;U��؉E�uhd�j j8h�)j�Ŏ������u̃}� u0�x����    j j8h�)h�)hd��{������   ��  �U� 3��} ����#E��;E��ىM�uhH)j j=h�)j�M�������u̃}� u0� ���� "   j j=h�)h�)hH)�������"   �J  3��} ���E�}� uh$)j j>h�)j��������u̃}� u0蚭���    j j>h�)h�)h$)蝥�����   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R��������P�E��P�MQ������3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V������M��UR�F�������蹫���0^]������������������������̋�U��Q�E�    �	�E����E��}�-s�M��U;��u�E�����7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]��������������������������������������������̋�U��Q�����E��}� u	�   ���ڪ���M�3���]�������������������̋�U��Q3��} ���E��}� u!h �j h�   h�*j�Ŋ������u̃}� u%j h�   h�*h`*h �胢�����   ��S����U� �3���]������������������������������������������̋�U��Q�����E��}� u	�   ��� ����M�3���]�������������������̋�U��Q3��} ���E��}� u!h �j h�   h�*j��������u̃}� u%j h�   h�*h�*h �裡�����   �虒���U� �3���]������������������������������������������̋�U��Q�.����E��}� u	������E�����]���������̋�U��Q������E��}� u	������E�����]���������̋�U���,���3ŉE��EP�M�Q�m������U�Rj j���ċMԉ�U؉Pf�M�f�H��������U�B�E�M��U��E�Pj j(h�+h�+h+�M�Q�UR�EP詩����P�X������M�U�Q�E�M�3��˫����]���������������������������������������������������̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]���������������������������������������������������������������������������������������������̋�U����X��E��M�����Ƀ��M�uh�,j j*hX,j�N�������u̃}� u+�����    j j*hX,h(,h�,�������E���E�X��E���]��������������������������������̋�U��X�]����̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�.j jh .j萅������u̃}� u0�C����    j jh .h�-h�.�F������   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U�E�Ph�   �M��Q�х����3҃} �U��}� uh�-j jh .j�˄������u̃}� u0�~����    j jh .h�-h�-聜�����   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U��E�Ph�   �M��Q�̈́������-��t3�t	�E�   ��E�    �M܉M�}� uh<-j jh .j调������u̃}� u-�c���� "   j jh .h�-h<-�f������"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9<�s
�<��E���M+M����U+щU؋E�Ph�   �M+M��U�D
P������3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ����������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����������������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U��W�}3�������ك��E���8t3�����_��������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��������������������������������������̋�U��j襙����]���������������̋�U��3�]�������̋�U����E���]��E���]���������̋�U����E�    �E�    �	�E����E��}�$}Z�M��<���uK�U�k���`��E������M����M�h�  �U�����P�D"��u�M�����    3��뗸   ��]��������������������������������������̋�U����E�    �	�E����E��}�$}O�M��<��� t@�U��<���t3�E������M��U�R�P"j�E�P�9������M�����    ��E�    �	�U����U��}�$}3�E��<��� t$�M��<���u�U������E�M�Q�P"뾋�]��������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�   �=�� u�����j�������h�   �܀�����E�<��� t
�   �   h  h�.jj�v�����E�}� u�s����    3��   j
�F~�����E�    �M�<��� uDh�  �U�R�D"��u"j�E�P�Ï�����"����    �E�    ��M�U�����j�E�P蒏�����E������   �j
跎����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��E�<��� u�MQ��v������u
j��������U����P��"]�����������������̋�U��E����Q��"]��������̋�U��EPj ��"h�   �����]����������������̋�U��j�h��h)d�    P�ĘSVW���1E�3�P�E�d�    �} u3��   j�v������u3��oj�[|�����E�    �EP�MQ��蠘���URj �EP�MQ�UR�M�觙���M��{����E���J����E������   �j������ËE�M�d�    Y_^[��]��������������������������������������������������������������̋�U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� �����������������̋�U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]�������������������̋�U��j�h��h)d�    P�ĘSVW���1E�3�P�E�d�    �} u3��   j�Et������u3��pj�z�����E�    �EP�MQ��������U R�EP�MQ�UR�EP�M������M�躘���E��艊���E������   �j�(�����ËE�M�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�M��M�茗���M���,聗���E�4��4��0��} t�U�<��E�8���8�    �<�    �M���,�(��U��$��E�@��M�D��H� �E���]� ��������������������������������������������̋�U���H�M��M���{���M��{���=4� ��   �4����?uG�4��B��@u8�0����0��U�R�����Phl7�E�P�a�����P�M��Cp���v�4����?uS�4��H��$uEj �U�R� �����P�M��p���M��rw����u�4��0��M�Q�9����P�M���o����U�R�"����P�M���o���M��/w����u	3��  �?�M��w����t�ώ����u�0����t�4�R�M��s�����E�P�M��vo���=8� u2�M�詔�����<�jh��<�Q�Z������E��U��8��=8� ��   �<�P�8�Q�M��L����8��U�E�E�M����tY�E���� u0�U���U�E��  �M���M�U���� u�M���M�����U�E��
�U���U�E���E�띋M�U���8���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M�jPhX��M������X���]���������������̋�U���h�L�����tH�@�%�����@�j �M�Q�n�����@���    �@��E�P�M�~����E�  �  �0����?�t  �0����0��0����?uK�0��H��?u=�U�R�{|�����0����t�0����0���E�P�M�����E�9  �M�Q�_y�����M��Jt���E�M��{���E��M�������u�U�R�M迃���E��  �0������   �0����@��   �M�Q诗�����M��9�������   �H���tn�H� �E�P�M�Q�M��q��P�M��Ql���0����@t>�M�Q�Z�����P�M��.l���U�R�E�Pht7�M�Q�M��&~�����Tq��P�M��l���)�U�R�E�Pht7�M�Q�M���}�����)q��P�M���k���}� t�M��.����}� t�M��x���M��k����u�M�������t�U�R�M藂���E��   �   �0����t�0����@ut�0����t�0����0�耊����t:�}� u4�M��$z����u(�M��Nv��P�M�Q衑�����U�R�M�����E�U��E�P�MQ�~������E�>�j�M�0����E�-�+�0����tj�M�����E��j�M�����E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��0����?uJ�0��B��$uj�MQ览�����E�;�$�0����0�j j �EP�6������E��j j�MQ�7�����E]�������������������������������̋�U���h���3ŉE�0����0�M�x5�}�	/�0����0��E�P�MQ�(��jl���E�;  �6  �M��t���0����?ubj �M�Q�ˇ����P�M���h���0���0����0���@t)�0����0��0������ك�Q�M��!l���  jh�7�0�R���  ����u�E�7�0����0��9jh�7�0�Q�ί  ����u�E��7�0����0���E�    �}� ��   �E�P�Β�����gy����twj�M�Q�M��+����U�R�ɍ����P�D����EЃ}� t�E�P�M��x���:h|7�M��x��hx7�M�Q�U�R�E�P�M�Q趂�������y��P�M��]n���:h|7�M��qx��hx7�U�R�E�P�M�Q�U�R�z��������oy��P�M��!n���N�E��t.�0����@u �M��Mr��P�M��,g���0����0��j@h0��M��ł��P�M��g���M��t�(��ci����u�U�R�(��f���E�P�M��}���E�M�3��ݐ����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �M��q���M��
q���E�    �E�    �0��������0����0����������������_�o  �������\��$�@��0����0�j�M����E�  �M��p���M����   �U�R裎����Pj<�E�P�4v����P�M��l���M������ȃ�>u
j �M��x���j>�M��n����} t�U��0����u�U�R�M��{���E�  �0����0��0��M�j j �U�R�z����P�M���d���Eܣ0��M��ix����u*�0��Q���1u�E�Pj~�M�Q�wu����P�M��d���M��3x����u�U�R�M��:k���E�P�M�_{���E�v  �%  �0��Q��� 5P�M��*u���  �E�   �0��Q����4P�M��u����  �0��������0����0����������������_��  ����������$����0����0�j�M��}���E��  �0��B����5Q�M��{t���F  �0��B����5Q�M�d���E�  �  �0��B����5Q�M���c���M��'p���U�R�M�/z���E�F  ��  jh�3�E�P�-d�����M��t���M�Q�M��y���E�  �0��B���t5Q�M�c���E��  �0��B���t5Q�M��s��j j �U�R�H�����P�M��b���M��Nv����u�M��l����tj�M�|���E�  �E�P�MQ�M��g���E�{  �  �  �0��B���t5Q�M��*s���0����uj�MQ�M��ϊ���E�4  �0����0�E�x�}�rj�M�2|���E�  �M���7R�M���r���0��������0����0������������������0�����������>  ������$�P�j �E�P��a�����M�Q�UR�E�P��t���Qj ��|���R�M��e�����f�����f���E�^  �  �E�P�M�Q�M��sf��j,��d���R��l���P�ԋ��������d��P�M���g��j,��T���Q��\���R謋�������d��P�M��g��j,��D���P��L���Q脋�������~d��P�M��g��j)��4���Rj ��<���P��x�������Td��P�M��Wg��j'�MQ�M��=d���E�  �;�U�R�EP�M��e���E�w  �!�0����0�j�M�{z���E�T  ��  �0��B���t5Q�M��q����  �0���� ����0����0��� ��������������� t������0t!�N�0����0�j�M��y���E��  j h�7�M�Q�`�����M��Dq���U�R�M�v���E�  j�M�y���E�  �0  �0���������0����0���������������������A������������	��   ��������l��$�d��0��Q����5P�M�_���E�  �0��Q����5P�M��_���0����?u5��,���P�n����P�M��e���0����@u�0����0����$���Q��j����P�M��Me��h�7�M��}���U�R�M�eu���E��j�M�x���E�n�j�M�x���E�]�j�M�px���E�L�}� t
�M��t���-�M���q����u!�E�Ph�4�����Q�y����P�M���]���U�R�M��t���E��]ÍI ����ȼ����� V�w�����	�'���I�þȾ������ 	

����������'�        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M���Z���0���0����0���@u�0���0����0���_tj�M�4t���E�   �0����0�j �U�R�r����j �E�P�r�����0����t�0����@t�0����0��ա0����u�0����0�j�M�s���E��0����0��M�Q�M�Up���E��]��������������������������������������������������������������������̋�U����   �M��d���E� �M��Z`������  �0������  �0����@��  �H���t�I���u�E�P�M�o���E�(  �M��Gl����uE�M�Qht7�U�R�s����P�M��pX���E���t�M�Qj[�U�R�>i����P�M��MX���E� �0����?�  �0����0��0����@�����@�����$��@�����@���%��  ��@��������$����0��B��_ua�0��Q��?uR�0����0��M�Q�U�Rj j �E�P�F���������\��P�M��W���0����@u�0����0��@�M�Q�U�Rj'�E�P�M�Q�f����Pj`�U�R�:h�������[�����\��P�M��;W����   �0����0��M�Q�U�Rj j�E�P��l�������P\��P�M��W����   j@h0��M��r���M�Qh�7�U�R��q����P�M���V���(��5Y����u�E�P�(��aV���w�0����0��U�R��|���Pj]�M�Qj j�U�R�5l�������8Z�����[��P�M��hV���E��*�E�P��l���Q��t���R�U~�������[��P�M��8V���.�E�P��\���Qj j��d���R��k�������W[��P�M��V�������0����<�����<��� t��<���@tW�W�M��i����tj�M��ZY���;�U�R��D���Pht7��L���Qj��T�����o�����g������Z��P�M��U����
j�M��Y���U�R�M�rl���E��]Ð��!�2�n��� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����0����uj�M�Zn���E�T�R�0����?u3�0����0�j �U�R�(l����Pj-�EP��d�����E��j �MQ�l�����E��]�������������������������������������̋�U���   V�E�    �0����Qu�E��7�0����0��0����uj�M�m���E�S  �N  �0����0��   �0����9��   �}� tG�0�� ��/��E��U��0����0��U�R�E�P�M��p��P�M�Q�U�R��m�����E��4�0�� ��/��E��U��0����0��U�R�E�P�M��>p���E��M��M�U�R�M�i���E�  �  �E�    �E�    �0����@��   �0����uj�M�l���E�L  �W�0����A|7�0����P*�E��U���W���ȋ�0����A���M��u��j�M�,l���E��   �0����0��e����0���0����0���@tj�M��k���E�   �M��tX�}� t&�U�R�E�P�M��o��P�M�Q�U�R�l�����E���E�P�M�Q�M���n���E��U��UЋE�P�M�Nh���E�V�T�}� t&�M�Q�U�R�M���n��P�E�P�M�Q�8l�����E���U�R�E�P�M��n���E��M��M��U�R�M��g���E^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����0����u3���   ��   �0����0|8�0����9*�0����/�M��0����0��E��   �   �E�    �0����@tY�0����u3��k�7�0����A|$�0����P�U����0���T
��U������2�0����0�뚋0���0����0���@t�����E���]����������������������������������������������������������������������̋�U����   �0����?u�0��B��$tj�M�i���E�  �0����0��$��U��(��E̋,��M���\����t���M��t���M��t����\����$��E��(��MЉ,��M��sY���M��kY���E� �0����?u/�0����0��U�Rj��T���P�v����P�M��N���jj��L���Q�c����P�M���M���M��a����t�H��U���up��D���P�w����Pj<��<���Q�^����P�M��}T���M��n���Ѓ�>u
j �M���v��j>�M���v���E��t�0����t�0����0��M��$��Ủ(��E��,��M�Q�M�Bd���E��]�����������������������������������������������������������������������������������������������������������������̋�U���|���3ŉE��E�   �M���W���I��M��	T�����  �0�����  �0����@��  �}� t	�E�    �
j,�M��u���0����0�U�x4�}�	.�0����0��M�Q�U�R�,��zO��P�M���R���  �0��E�M��W���0����Xu�0����0�h8�M���\���%  �0����$u7�0��H��$t)�0����0��E�P��s����P�M��K����   �0����?��   �E�P�4v������\����tkj�M�Q�M��h���U�R�/q����P�D����Eă}� t�E�P�M��"\���.hx7�M�Q�U�Rh�7�E�P�(f�������]��P�M��K���.hx7�M�Q�U�Rh�7�E�P��e��������\��P�M���J����M���U��P�M�Q�O����P�M��J���0�+U��~�,��M����u�E�P�,��7J���M�Q�M��GQ��������I� �U�R�M�`a���E�M�3��mt����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE�0���M��0����0��E�������������R��  �����������$�p��EP�t�����E�  �0����@u$�0����0�h8�M��I���E�S  �3��D���Q�MX����P�URh�4��L����I�����)N���E�  �EP�X�����E�
  �M�Q�zs�����U�R�ns�����M��[������   �M��[����t{jd�E�P�M��e����uj�M�b���E�  �M��M��U���-u�E��E��E�.��E�.�M�Q�URje��4���P�M�Q��<�����H������K�����hM���E�]  �j�M�Ib���E�I  ��x���R�r�����OY����tSj��h���P��x����e����h���Q�m����P�D�����d�����d��� t��d���R�M�MH���E��  �E���Du5hx7�MQ��x���Rh�7��,���P�b�������xY���E�  �3hx7�MQ��x���Rh�7��$���P�Nb�������CY���E�m  �h  j j ��\���Q��\���������R��q������\���P�M��]���E�/  j{��T����c���M�������������H|3������J~�(�����R�V����P��T����sM��j,��T�����o���E���������������F������������wx�������$��������P�q����P��T����M��j,��T����o�������Q��p����P��T�����L��j,��T����jo��������R��p����P��T�����L��j}�EP��T����I���E�-�+�0����0�j�M�
`���E�j�M��_���E�M�3���o����]Ë�5�����V��B�1���S� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �M��O���i���E��M�<K���E��}���  uj�M��]���E�  �B�}���  u�EPj�MQ�Y�����E�  ��}���  u�UR�M�}Z���E�j  �E�% �  �0  �M��� �  t�U���   3���   ���������M��� `  ��Ƀ����������� t�U���   �� �����E�%   �� ����� ��� t>�M��� �  t�U���   3���   ���������
ǅ����    ������ ��
  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ t|�M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� @  tM�E����t/�5J����t&�U�R��O����Pj �E�P�R����P�M��A����M�Q��O����P�M��dc���U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t�E�%   ��������M���   ������������ �-  �U��� �  t�E�%   3�=   ���������
ǅ����    ������ ��   �U�R�-X����P��|���Pj{�M�Q�M�nD������E��P�M��jG���U�R�9L�����_����u1hH9��l���P�M�Qj,��t���R�PQ�������rR��P�M��$G��hD9�M���^���E�P��k�����D����tR�k����tI�T_����u@�M�Q��T���Rj ��\���P�M�Qj ��d���R��P�������C�����3E��P�M���?���  �M���J���M���J���M���J���M���J���M���J���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ �"  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t[�M���   ��   uJ��L���R��f����P�M���>����D���P��f����P�M���>����<���Q��f����P�M��>���k�U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t'�E�%   =   u��4���Q�af����P�M��<>����,���R�If����P�M��$>���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t8�U��� �  t�E�%   3�=   ���������
ǅ����   ������ u;�G����t��$���R�dT����P�M��==��������P�JT����P�M��_���A����tO�h����t,�M�Q�����R�����P�h�������6B��P�M���<��������Q�qh����P�M��^���������R�Wh����P�M��^���M�`P����uA�M��TP����u)��[����u �EPj ������Q�eM����P�M��@C����UR�M��f<���E�    �M��oG���}� tNj ������P� H����Ph@9������Q�@W����P�M���B���I[����t�U�R�M�
S���E��  �bj h�j�T���������������� t��������F���������
ǅ����    �������E��M�Q������R�jG����P�M��;���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ ��  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M���   ��   uzj,������R�E�P������Qj,������R�E�P������Qj,������R�E�Ph09������Q�U�������G>������?�����9>�����?�����+>��P�M��.A���   �U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� tB�E�%   =   u3j,������Q�U�Rh 9������P��T�������=��P�M��@���h9�M��oX��hH9������Q�M���K��P�M��y@��j)��x���R������P�ZY����Pj(������Q�kJ�������<=��P�M��?@���U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� ��   �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t:�M��� �  t�U���   3���   ���������
ǅ����   ������ u�M�Q�M��m?���K����t��p���R�H����P�M��L?�����h���P�H����P�M��NZ���Tc����t�}� t�M�Q�M��K8���U�R�M��?8���  �EP�M���>���M��� �  u.�U��� |  �� h  u�E�P�MQ�cR�����E��	  �1  �U��� �  u,�E�% |  = p  u�M�Q�UR�=<�����E�	  ��  �E�% �  u]�M��� |  �� `  uLhD9�UR��X���P�lJ����P��P���Qj{��`���R�M��2;�����<�����uI���E�N	  �  �E�% �  u.�M��� |  �� |  u�U�R�EP�H�����E�	  �[  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th�8�M��U���  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th�8�M��UT����   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tI�M��� �  t�U���   3���   ���������
ǅ����    ������ thp8�M��S���0�M��� �  u%�U��� |  �� x  u�E�P�M��K���E�  �M��� �  t�U���   3���   ����|�����M��� `  ��Ƀ���|�����|��� t�U���   ��x�����E�%   ��x�����x��� ��   �M��� �  t�U���   3���   ����t����
ǅt���    ��t��� u:�M��� �  t�U���   3���   ����p����
ǅp���    ��p��� t#�M�Qh@9��H���R��N����P�M��3����E�P��@���Q�JI����P�M��3���U��� �  t�E�%   3�=   ����l�����U��� `  ��҃���l�����l��� �x  �YY�����R  �E�% �  t�M���   3ҁ�   ��h�����E�% `  �������h�����h��� t[�M��� �  t�U���   3���   ����d����
ǅd���   ��d��� t!�M�Qhd8��8���R��M����P�M��2���E�% �  t�M���   ��   �s  �U��� �  t�E�%   3�=   ����`�����U��� `  ��҃���`�����`��� t�E�%   ��\�����M���   ��\�����\��� �$  �U��� �  t�E�%   3�=   ����X�����U��� `  ��҃���X�����X��� t�E�%   =   ��   �M��� �  t�U���   3���   ����T�����M��� `  ��Ƀ���T�����T��� t�U���   ��   tU�E�% �  t�M���   3ҁ�   ��P�����E�% `  �������P�����P��� t2�M���   ��   u!�U�RhX8��0���P�L����P�M���0����W�����  �M��� �  t�U���   3���   ����L�����M��� `  ��Ƀ���L�����L��� tl�U��� �  t�E�%�   3Ƀ�@����H�����U���   3���   ����H�����H��� t&�M�QhL8��(���R�\K����P�M��>0���Z  �E�% �  t�M���   3ҁ�   ��D�����E�% `  �������D�����D��� tp�M��� �  t�U����   3����   ����@�����M���   3ҁ�   ��@�����@��� t&�E�Ph<8�� ���Q�J����P�M��/���   �U��� �  t�E�%   3�=   ����<�����U��� `  ��҃���<�����<��� tb�E�% �  t�M����   ��Ƀ���8�����U���   ��҃���8�����8��� t!�E�Ph08�����Q��I����P�M���.���U��� �  t�E�%   3�=   ����4�����U��� `  ��҃���4�����4��� t�E�%   ��0�����M���   ��0�����0��� t*�M����u!�U�Rh$8�����P�gI����P�M��I.���M���   t!�U�Rh8�����P�;I����P�M��.���M�Q�M�E���E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���x�E�    �0����_u�U��� @  �U��0����0��0����A�  �0����Z�  �0����A�E��0����0��U��� �  �U��E���t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M�U����U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U��E��E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E܋M܉M��;�U��� �  t�E�%?����E���M��������M؋U؉U���E���  �E��k  �E����Eԃ}���   �M��$��	�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M̋ỦUЋEЉE����E���  �E��  �  �0����$��  �E� �0����0��0���Uȃ}�R�]  �E����	�$��	�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  �0��Q��Pu�0����0��0����0��0���Eă}�Q��   �M���T	�$�@	�0����0���J���  �0����0��0����0|C�0����95�0���0��D
ѣ0��J���E��M���   �M��E��-  ��E���  �7�0����0��UJ���	  �E���  �E���  �E���  �E���  ��  �E���  �0����0���  �E��0����0��0����0|�0����5~$�0����t	�E���  ��E���  �E��z  �0����0�E��M��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��M���t�U���    �U���E�%�����E��M����M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  �0����0���  �0����0��  �0����8��  �0���U�0����0��M�������M��U�U��E���0�E��}��?  �M��$��	�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C�0����9u�0����0��E���  ��0����t	�E���  ��E���  �E���]ÍI ����|���j���S�����'�>�U���j������� 																																																																					��������� �����J 	� 	� 	� 		'	9	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j �S&����P�M��L���0����tl�0���E�0����0��U�U�}�0t�}�2t�}�5t(�5h8�M���9���&�E�P�0����P�M��	"���j�M�l5���E�(�
j�M����hL9�M��9���M�Q�M�2���E��]���������������������������������������������������̋�U���@�M���%��j j�E�P�c0����P�M�����M��"����uN�0����tA�0����@t4�U�R�E�Pht7�M�Q�U�R�E�������k,�������P�M��J���0����@u�0����0��b�0����tj�M�����J�M���-����tj�M�����2�U�R�E�Pht7�M�Qj�M��4������+�������P�M������U�R�M�0���E��]��������������������������������������������������������������������������̋�U����0�����  �0����A�E��0����0��}���   j�M��^3���������   �U�����U��}���   �E���		�$��	j�#����P�M���)���|j�{#����P�M��)���gj�f#����P�M��)���Rj�Q#����P�M��)���=j�<#����P�M��z)���(j�'#����P�M��e)���j�#����P�M��P)���U�R�M�R/���E� �j�M�2���E��j�M�n2���E��]ÍI +	@	U	j		�	�	�	 ��������������������������������������������������������������������������������������������̋�U��0����@u"�0����0��EP�M��-���E���MQ�UR�������E]�����������������������̋�U��� �EP�M��-���0���U��}� t�}�?tq�}�Xt��   �E�Pj�MQ��,�����E��   �0����0��M��*����th8�M�o���E�   ��E�PhP9�MQ�1�����E�w�0����0��E�+�j �M��!��P�E�P�M�Q�U�R��?����P�M��c���E�P�MQ������E�$�U�R�M�?-���E��E�P�MQ�r�����E��]�������������������������������������������������������������������������̋�U���<�M��� ���0���Mȃ}�B��  �U���	�$� 	�MQj�UR�+�����E�j  hl9�M��o&���M�-)����u
j �M��>���EP�M��[,���0����0��E��4�U�R�M��Y*��P�E�P�MQ�������E�   �0��B��$t<�0��Q��u�EPj�MQ��*�����E��  �j�M�/���E�  �0����0��0���Mă}�T�o  �U���|	�$�X	�0����0��UR�EP�I9�����E�Y  �0����0�j�UR�EP�������E�0  �0����0��E�+�j �M��K��P�U�R�EP�M�Q�=����P�UR�.�����E��   ��   hl9�M���$���M�'����u
j �M��0=���EP�M���*���0����0��E�|4�U�R�M���(��P�E�P�MQ�A�����E�z�0����0�j�M�-���E�\�G�0����0�hX9�M����E�;�&�MQj�UR�K)�����E�"j�M�v-���E��EP�MQ�(-�����E��]Ë�v	�	�	�	�	 ��	z	�	�	<		�	�	�	 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �0���M�}�XtD�}�Zt�`�0����0������t	�E�0��E�9�E�P�M����E��   �0����0�h8�M����E��   �U�R��;�����M��5������   �0���M�}� t�}�@t`�}�Zt�v�U�R�M�'���E�   �0����0�������t	�E��9��E�x9�M�Q�U�R�M��j"��P�M�M'���E�>�0����0��M�Q�M�/'���E� j�M�^*���E���U�R�M�'���E��]��������������������������������������������������������������������������������������������̋�U���,�E�   �M�����M��������  �0����@��   �0����Z��   �}� t	�E�    �
j,�M��8���0������   �0����0�M�x3�}�	-�0����0��E�P�M�Q�$��X��P�M������k�0��U�M�����P�E�P������0�+M��~�$��0����u�U�R�$��\���E�P�M��l���0�;M�u
j�M�����j�M�����������U�R�M�i%���E��]����������������������������������������������������������������������������������������̋�U���(�0����tg�0����Zu'�0����0��M�����P�M��$���E�^�0j)�UR�E�P�w-����Ph�9�M�Q�(�������Y���E�,�*j)�URj�E�Ph�9�M��#�����!6�����+���E��]�������������������������������������������������������̋�U���x�0�����k  �0���E��0����0��E� �E������M�� ���U��U��E���C�E��}��   �M����	�$��	hp:�M�����?  hh:�M�����-  hd:�M��{���  h\:�M��i���	  hT:�M��W����  hL:�M��E��hD:�M���*����  �E����E���  �0���U��E�E��0����0��U��U��}�Y�8  �E���	�$��	�E������(  h<:�M������  h4:�M�����  h(:�M������   h:�M������   h:�M������   h:�M��o���   h�9�M��]���   h�9�M��K���   �0����0��E�P�����P�M��3���M�������t�M�Q�M�"���E�~  �R�UR�E�P�%����Ph�9�MQ�&�����E�R  �0����0�j�M��\���h�9�M�����Qh8�M�����B�0����0��M�Q�s����P�M��
���M��9����t�U�R�M�q!���E��  �}����   �E��E��M���C�M��}���   �U���x	�$�h	�M�Qh�9�U�R�7%����P�M��
���e�E�Ph�9�M�Q�%����P�M���	���E�U�U��E���E�E��}�w/�M����	�$��	�E�Ph�9�M�Q��$����P�M��	���M�_����u�URj �E�P�|����P�M��W���M�Q�M�| ���E��   ��   �M�����UR�M��[ ���}��uF�M��m2���E�P�M�Q�U�R�������M�������uh�4�M���'���E�P�M� ���E�}�M�����tA�M���t$h�9�M������U���th�9�M��'����E���thl9�M�����M�Q�U�R�EP�������E���MQj�UR������E��]�`	r	�	�	�	�	�	�	`	�	o	   










	�I 6		H	Z	l	~	�	6	*	�	�	�	Q	 	
��	�	&	k	 �I M	k	     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�$����t�%����u	�E�   ��E�    �EЉE��M������0���U̡0����0��M̉Mȃ}�Y��   �U����	�$�t	�0����0�h�:�M����E�   h�:�M��I���kh�:�M��:���\h�:�M��+���Mh�:�M�����>h�:�M�����/��#���E��U�R�+����Phx:�E�P� ����P�M������M������}� t�M�Q�M������U�R�6����P�M�����E�P�M����E��]Ë��	�	�	�		�	�	0	 ���������������������������������������������������������������������������������������������������������������������������������̋�U��EP�������E]����������̋�U����M�����0������   �0���E�M��0�M�}�wH�U��$��	h�:�M��*���>h�:�M�����/�-h�:�M��
���hL:�M������j�M�;���E�~�0���M�0����0��E�E�M��1�M�}�w/�U����	�$��	�M�Qh�9�U�R�����P�M�����E�P�M����E��j�M����E��]��	�	�	�	�	�			b	�	    ��������������������������������������������������������������������������������������������̋�U����   �0����u�URj�EP�������E�  �0����6|�0����9~ �0����_tj�M�����E��  �0����6�U��0����0��}�)u[�0����t2�0����=�M��0����0��}�|�}�~�E�������EPj�MQ������E�M  ��}� |�}�~�E������}��uj�M����E�   �M������UR�M������E����  �M�Qht7�U�R�����P�M�� ���0����t5�U�R�E�P�M�Q�+����Pj �U�R�T���������P�M��\ ����E�Pj�M�Q�I����P�M��? ���0����t1�0����@u�0����0��j�M�F���E�J  ��M�Qj�UR�������E�.  �	����t�E�P������P�M��������M�Q������P�M��!���U���tS�����t5�E�P�M�Q�U�R������Pj �E�P�f���������P�M��n�����M�Q�����P�M��?!���5����t)�U�R��x���P�M�Q��*�������v��P�M��'������p���R�*����P�M��� ���M�����u.j)��`���P�M�Qj(��h���R�����������P�M������j h�j��������\�����\��� t��\�����	����0����
ǅ0���    ��0����E��M�Q�U�R�=
����j)��D���P��T���Q�*����Pj(��L���R�;���������P�M����������t�E���t�M�Q�M����������t��<���R�$����P�M��������4���P�
����P�M������}� t�M�Q�M�������j�M����E��U�R�M����E��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����0������   �0����6|�0����9~�0����_un�UR�M�������M������u$�M������u�M�}����u�EP�M������M������u�MQ�M������U�R�EP� �����E�   �>j �MQ�UR�EP�M�Q�g%�����U�3Ƀ�*��Q�U�R�EP�8������E�m�kj�M������MQ�M��=���M�E����u�UR�M��L���M�-����u"�M�!����u
j �M��$���EP�M�����M�Q�M�C���E��]��������������������������������������������������������������������������������������������������̋�U���4�M������0����0��0���UЀ}�At�}�BtN�}�C��   �   �} u%�E����&u	�E̤4��Ē4�E�M̉�0����0��  �} tj�M����E�}  �E� j>�M��(���0����0��N  �U��4�0����0��3  �0����t�0��H��uj�M����E�  �} tj�M����E��   �0����0���0��Q�DЉE�0����0��}�v/j,�M��v���U�3�PR�M����P�M�Q�M�����P�M��\���j>�U�R�M�����P�M��E����0����$u�0����0��j^�E�P�M������P�M������0����t�0����0��
j�M������M��y ���M�Q�M�����E��M�����E��]�����������������������������������������������������������������������������������������������������������������������������������������������������̋�U���$  �M��2���E� �0�����  �0����$u8�MQ�U�R�EP�M�Q�S�����M������u�U�R�M�����E�  �0���0��3҃�A����+��+ʉM�M�����M�����E�   �E艅����������t������tw��������   �  �3�����tW�v����tN�M���
����u/j������P�M�Qj �U�R�M���������$	��P�M��
����j�����P�M������   �������tN�M��
����u/j
�y����P�E�Pj �M�Q�M��~���������P�M������j
�J����P�M�����`�u�����tN�M��;
����u/j	� ����P�U�Rj �E�P�M��%������o��P�M��U����j	�� ����P�M��/����E�    �}� t|�0����0��0����$u8�MQ�U�R�EP�M�Q�o�����M��	����u�U�R�M�����E�  �0���0��3҃�A����+��+ʉM�}� �)����0����t�0����0��}���  �EP�M��$����M�Q�U�R�M�����P�M��a����M��	����u)�E�P��|���Qj �U�R�M���������{���P�M��,����M�������u,�E�P��l���Qj ��t���R�M���������C���P�M�������E���  �} tj�M����E�  �M���tz�E�Pht7��d���Q������P�M������0����t,�M�Q��T���R��\���P�����������P�M��n�����M�Qj��L���R�X
����P�M��N����$�0����t��D���R�T����P�M�����0����uj�M������/�0���0����0���@tj�M�$���E�  ������t[�U��������������t�B�} tj�M�����E�t  �E�P��4���Q��<���R�������������P�M������#�E����u��,���Q�����P�M��B���U��t!�E�Ph�:��$���Q�O����P�M��1����U��t!�E�Ph�:�����Q�&����P�M������} ��   �M�������   �M�3
����u�M�����t:�M�w����t�UR�M�������EPj �����Q�����P�M��j����@�UR������Pj �����Q�URj �����P�[�������,���������P�M��(����*�M�����u�MQj ������R�!����P�M�������M��E���E���t�M��M���M�Q�M�		���E��   �j�M�3���E�   �   �} ux�M�����ul�M�	����u�M�z����t�URj�EP������E�u�9�MQ�URj ������P�MQj������R��������;����������E�:�8�} u%�M�����u�EPj�MQ�J�����E��j�M�s���E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����0�����  �} t]�0����XuO�0����0��M������th8�M������E��   ��URhP9�EP�
�����E��   �0����Yu%�0����0��MQ�UR�������E�   �EP�M�Q������M�Y�����t �U�Rh;�E�P�	����P�M������*�M�����t�M�Qh�:�U�R�w	����P�M��Y����E�P�M�J���E���MQj�UR�5�����E��]��������������������������������������������������������������������������������̋�U���   �0�����s  ������E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M��V
�����9�����C���P�MQ�x�����E�  �  �M��y����M�����th�4�M������M��2 ����tR�U��E����E���tB�0����t5j]�E�Pj �M�Q�F����Pj[�U�R�������������P�M�����뢋M� ����u^�M�����t�E�P�M�Q�M����P�M������7�U�R�E�Pj)�M�Q�URj(�E�P���������P����������P�M������M�Q�U�R�������M�����E�P�M�Y���E�   �   �M�������uSj]��|���Qj�U�Rh;�E�P�MQj(�U�R���������#���������������P�EP�������E�?�=j]��d���Qj��l���Rj[��t���������y��������P�EP������E��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j'�EPj �M�Q�<����Pj`�U�R��������������E��]�����������������������̋�U����E�+�j�M������P�E�P�M�����P�MQ�-�����E��]����������������������̋�U��Q�E��4�E�P�MQ�UR�EP������E��]��������������������̋�U��Q�E�+��E�P�MQ�UR�EP�� �����E��]��������������������̋�U��EP�MQ�UR�EP� �����E]��������������̋�U��j�EP�������E]��������̋�U��j �EP�������E]��������̋�U��j �EP������E]��������̋�U��EP�MQ������E]������̋�U��Q�0���M��}� t)�}�At�0�0����0�h;�M�����E�j�M�?���E�j�M�0���E��]���������������������������������̋�U���@�EP�M������M��������b  �0�����Q  �E�P�M�Qj �U�R�E�P����������7���������P�M��g����M��Q������  �0����@��   h(;�M������M��"�������   �0������   �0����@txj'�M�Q�U�R�����Pj`�E�P�������������P�M������0����@u�0����0��M�������t�0����@th$;�M��<���Z����M��|�����t �0����u
j�M�����j}�M�����0����@u�0����0��'�M��1�����t�U�Rj�E�P�*�����P�M�� ����M�Q�M�����E��]����������������������������������������������������������������������������������������������������������������̋�U��EP�W������E]����������̋�U����E�+�j �M��|���P�E�P�M��o���P�MQ�������E��]����������������������̋�U����EP�M�����h(;�M�����M�Q�#����P�M������j}�M��<���0����@u�0����0��U�R�M������E��]��������������������������������̋�U���,j h�j�������E��}� t�M������E���E�    �EԉE�M�Q�U�R��������EP�M�Qj �U�R�E�P�y���������������o���P�M�� ����M�Q�M�����E��]������������������������������������������������̋�U��@��������]����������̋�U��@�%   �����]��������̋�U��@��������]����������̋�U��@��������]����������̋�U��@��������]����������̋�U��@���`3Ƀ�`����]�������̋�U��@�%�   �����]��������̋�U��@�%   �����]��������̋�U��@�%   �����]��������̋�U��@�%   ]���������������̋�U��@�%    ]���������������̋�U��@�% @  ]���������������̋�U��@�% �  �����]��������̋�U��@�%   �����]��������̋�U���������t�E���5���M���5��]���������������������̋�U��@��������]����������̋�U��EP�MQ������]�������̋�U����M�E������E�} t�MQ�U��Ѓ���   ��   �} w�E   �M�Q;U��   �}   v3��   jh�h  �;������E��}� t�M�����E���E�    �E��E��}� tA�M�y t�U�B�M���U�E��B��M�U��Q�E�M��H�   +U�E�P�3��!��M�Q+U�E�P�M�Q�E�H�D
��]� ���������������������������������������������������������������������̋�U��Q�M��E��     �E���]�������̋�U����EP�MQ�UR�M���������O����E��]���������������������̋�U����EP�MQ�UR�M������������E��]����������������������̋�U����EP�MQ�UR�M��;�����������E��]����������������������̋�U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]�����������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��Z����E���]� ������������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��} tdj h�j�.������E��}� t�EP�M��?����E���E�    �M��U��E����Ƀ�������   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ���������������������������������������������������������������������������������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ��"  ���E��}� v�U�R�EP�M������E���]� ���������������������������������������������������������������������̋�U���V�M�E�H�� ����U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E��     �M�Q�������E�P�M�Q�������E�P�M�Q�������E�P�M�Q������E�P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	������t�U����U���E�H�� ������U�J�   ������E�P�M�Q�M������U����t<�U�E���M�	���u�;�t�U�B% ������M�A�U��    �!�M�������u�E�H�� ������U�J��E�H�� ������U�J��E�H�� ������U�J�E�^��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��@�%   ]���������������̋�U���$���3ŉE��M܍E��E��M܋Q�� ����E܉P�M��    �U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%����M܉A�U�� �E����E�j j
�MQ�UR�������0�� �M��j j
�UR�EP�����E�U�MMu��U��E�+й   +�Q�U�R�M������E܋M�3��� ����]� ����������������������������������������������������������������������������������������̋�U���(���3ŉE��M؍E��E܋M؋Q�� ����E؉P�M��    �U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%����M؉A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U܃��U�j j
�EP�MQ�0�����0�� �U܈j j
�EP�MQ�H����E�U�UUu��E��t�M܃��M܋U��-�E܍M�+��   +�R�E�P�M������E؋M�3�������]� ��������������������������������������������������������������������������������������������������������̋�U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�\������M���U��: u�E��H�� ������U��J�E���]� �����������������������������������������������������������������������̋�U��Q�M��E��H����3�������]���������������̋�U��Q�M��E�3Ƀ8 ������]������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J�E���]��������������̋�U��Q�M��E��@������]�������̋�U����M��M�������u�E��H��	��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��M��������u�E��H��   �U��J��]���������������������̋�U����M��M�������u�E��H��
��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��    �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� @  �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� �  �U��J��]�����������������̋�U��Q�M��M�������t3���E���U����ȋ�Ћ�]�����������������̋�U��Q�M��M��a�����t2���E���U����ȋB�Ћ�]����������������̋�U����M�M�������uX�} u*�M��������Ej h��EP�R������E��M��M�} t �U�E�L�Q�UR�M������E��E��  ��} t�M� �E��]� �������������������������������������������̋�U��Q�M��M��q�����t�E��EP�MQ�U���M��	��B�Ћ�]� ����������������������̋�U����M�E�P�M��c����MQ�M������U�R�M�J����E��]� ����������������������̋�U����M�E�P�M������MQ�M������U�R�M������E��]� �����������������������̋�U����M�E�P�M�������MQ�M������U�R�M�����E��]� �����������������������̋�U����M�E�P�M��s����MQ�M������U�R�M�[����E��]� �����������������������̋�U����M�E�P�M��#����MQ�M������U�R�M�����E��]� �����������������������̋�U����M��} t_j h�j��������E��}� t�EP�M��R�M��h����E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ������������������������������������̋�U����M��M�������tb�E��tZ�M��������t�MQ�M�������?j h�j�������E��}� t�UR�M������E���E�    �E�P�M��H����E���]� ���������������������������������������������̋�U����M��M��l�����tu�} to�E���te�M�������t�UR�M��=����Kj h�j�N������E��}� t�EP�  ��P�MQ�M������E���E�    �U�R�M������E���]� ������������������������������������������̋�U��Q�M��M�������tG�M�e�����t�M����P�M��9����(�M��F�����t�EP�M�������M�R�M�������E���]� ��������������������������̋�U����M��M��,�������   �} ��   �M��������t�EP�M�������j�M�r�����t�M�f�����u@j h�j��������E��}� t�MQ�M������E���E�    �U�R�M��;�����M����P�M��B����E���]� ���������������������������������������������̋�U��Q�M��M��N�����tC�M�������u�}t�}u�EP�M��������} u��MQ�������P�M������E���]� ������������������������������̋�U����M��M��F�����t3�M������u'�M�-����E��E�%�   �M��Q�� ���ЋE��P�E���]� ���������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��Z����E���]� ������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�  ��P�UR�M��G����E���]� ���������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h�j�s������E��}� t�MQ�M������E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������̋�U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ�������U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ������������������������������������������������������������������̋�U����M�E�8 tj�M�������  �} ��   �} ��   �M�M��}� t�}�t�u�U�B% ������M�A�   j h�j�������E��}� t�U�P�M������E���E�    �M�U��E�8 u�M�Q�� ������E�P�[j h�j�������E��}� t�MQ�UR�M������E���E�    �E�M��U�: u�E�H�� ������U�J��E�H�� ������U�J��]� ����������������������������������������������������������������������������������������̋�U��Q�M��E�3Ƀ8	������]������̋�U��Q�M��E�� �����E���]�������̋�U����M�M��������uf�M�3�����uZj h�j�|������E��}� t�EP�M��Q����E���E�    �M��M��}� t�U����M��U��M�U��T��E��]� �����������������������������������������̋�U��Q�M��} |�}	~j�M�	����E�;�9�E��8�t
�M��U;~j�M������E���E�M��T�R�M�����E��]� ��������������������������̋�U��Q�M��E�� 0;�E���]�������̋�U��Q�M��M�������E�� @;�M��U�Q�E���]� �������������������̋�U��Q�M��   ��]��������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E;Es�M�U��B��M���M�E��]� �����������������̋�U����M��M��6����E�� P;�} tP�} tJj h��MQ�e������E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ�S  ����U��B    �E��@    �E���]� ������������������������������������������������̋�U��Q�M��E��@��]�������������̋�U����M��E��x t�M��Q�E��H�T
��U���E� �E���]����������������������������̋�U��Q�M��E��HQ�U��BP�MQ�UR��������]� ������������������̋�U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�"  ���EE��]���������������������̋�U����M��M��v����E�� `;�} t#�M������t�M������u	�E�    ��M�M��U��E��B�E���]� ����������������������������������̋�U����M��E��x t�M��I�r����E���E�    �E���]��������������̋�U����M��E��x t�M��I������E���E� �E���]�����������������̋�U����M��E��x t�MQ�UR�E��H�A����E���M�M��E���]� ��������������������̋�U��Q�M��M��(����E�� p;�M��U�Q�E��H����Ƀ�����U��J�E���]� ��������������������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E��x��,"�;��]�����������������̋�U��Q�M��E��xujh�;�MQ�UR��������E��]� ���������������������������̋�U��j�h�d�    P���3�P�E�d�    �����uM���������E�    j �������j����ۿ��j����Ͽ��j����ÿ���E������} |�}}�Ek��������M�d�    Y��]��������������������������������������������������������̋�U��Q�M��M��H����E�� �;�M��U�Q�E��M�H�U��B�����E���]� ����������������̋�U��QV�M��E��x }.�M��Q�E��H���Ћ��M��Q�E��H������M��q�U��B^��]��������������������̋�U����M��E��H�U��B��ȋB�ЈE��M���u�U��B�M��I��B�ЈE��E���]������������������������̋�U����M��EP�MQ�U��B�M��I��B�ЉE��M�;Ms�UR�E�P�M��Q�E��H��B�����E���]� ����������������������̋�U��Q�E�    �	�E���E�M���t�E����E���E���]����������������������������̋�U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]��������������������������̋�U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]������������������������̋�U��Q�E�    �}�wC�EP�������E��}� t�*�=�� u�T����    ��MQ�8�������u����UR�"������%����    3���}� u�����    �E���]���������������������������������������̋�U��Q�=�� u�����j� �����h�   ��������} t�E�E���E�   �M�Qj ���R��"��]�������������������������̋�U��QV�E�    �} u�4�EPj ���Q��"�E��}� u�$"P���������$����0^��]����������������������������������SVW�T$�D$�L$URPQQh0k	d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�x����   �C�&����d�    ��_^[ËL$�A   �   t3�D$�H3������U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�����3�3�3�3�3���U��SVWj Rh�k	Q�Y���_^[]�U�l$RQ�t$������]� ���������������������������������������������������������������������������������������������̋�U��E���]�����������������̋�U��Qj���������P��!�E��MQ��!���j��������E���]�����������������̋�U��} th<j jWh�;j���������u�j �q�����]���������������������������̋�U����P��!]�������������̋�U��Q���P��!�E��}� t�MQ�U�����u3���   ��]��������������������������̋�U��   ]����̋�U����    ]���������������̋�U���V3��} ���E�}� uh�<j jHhP<j���������u̃}� u-�����    j jHhP<h,<h�<������3��   �}�v�u����    3��~�} u�E   �URj ���P��"�E��MQ�URj���P��"�E��}� u:�}� @  w�M;M�w�x   ��t�U�U���$"P��������������0�E�^��]����������������������������������������������������������������������������̋�U����E�����j j�E�Pj ���Q��"��t�}�u	�E�   ��E�    �E���]�������������������������̋�U���V�E�E��} u�MQ苶������   �} u�UR�.�����3��   �E�    �}�w)�} u�E   �EP�MQj ���R��"�E���EP�����������    3��e�}� u	�=�� u%�}� t��$"P�������������0�E��1�MQ�d�������u�$"P����������R����03���J���^��]����������������������������������������������������������������������̋�U��Q�E�����j j ���P�0"��u�E������E���]�����������������̋�U������]����̋�U���<�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� uh�j jih(=j蒶������u̃}� u.�E����    j jih(=h=h��H���������  3Ƀ} ���M̃}� uh�<j jnh(=j�.�������u̃}� u.������    j jnh(=h=h�<�����������   �E�E��M��A����U��BB   �E�M�H�U�E��M�Qj �UR�E�P�������E��} u�E��Q�M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj �������EċE���]��������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ��������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�>�������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR���������]��������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR蒬������]������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�P�������]����������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�R�������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��������]��������������������̋�U��Q�E�E��M�Q�UR��������]����������������̋�U��Q�E�E��M�Q�UR�n�������]����������������̋�U��Q�E�E��M�Q�UR�EP�+�������]������������̋�U��Q�E�E��M�Q�UR�EP���������]������������̋�U��E��=   vh>j j8h�=j�>�������u̋UR�EPj ������]����������������������������̋�U����EP�M�豿���M����   vh>j jDh�=j�α������u̃}�|5�}�   ,�M������� ���   �U�Q#E�E�M��/����E��1�'�M��Ӱ������   �B�#E�E�M������E���M��������]��������������������������������������������������̋�U���(�EP�M��Ѿ���}�|6�}�   -�M��K�������   �E�B#M�M��M��{����E��   �M�����P�U�����   R蟲������t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M��ȯ��� �HQ�M�躯����BP�M�Q�U�R�E�Pj�M�螯��P�;����� ��u�E�    �M�������E���M�#M�M؍M������E؋�]������������������������������������������������������������������������������̋�U��=L� u�E����A#E��j �UR�EP�a�����]���������������������������U��WV�u�M�}�����;�v;���  ���   r�=` tWV����;�^_u�{�����   u������r)��$��y	�Ǻ   ��r����$��x	�$��y	��$�dy	��x	 y	Dy	#ъ��F�G�F���G������r���$��y	�I #ъ��F���G������r���$��y	�#ъ���������r���$��y	�I �y	�y	�y	�y	�y	�y	�y	�y	�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��y	���y	�y	�y	z	�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l{	�����$�{	�I �Ǻ   ��r��+��$�pz	�$�l{	��z	�z	�z	�F#шG��������r�����$�l{	�I �F#шG�F���G������r�����$�l{	��F#шG�F�G�F���G�������V�������$�l{	�I  {	({	0{	8{	@{	H{	P{	c{	�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l{	��|{	�{	�{	�{	�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]���������������������������������̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�������������������������������������������̋�U��j�h8�h)d�    P���SVW���1E�3�P�E�d�    �e��E�   �E�    �E�P谳������u�E�    �E������E��   �M+M�M܋U�R�E�P�֯�����E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]������������������������������������������������������������������������������̋�U��h"+��!���]���������̋�U��j�hX�h)d�    P���SVW���1E�3�P�E�d�    �e��׳���@x�E�}� t#�E�    �U��E�������   Ëe��E������E����M�d�    Y_^[��]��������������������������������̋�U��Q�f����@|�E��}� t�U��#�����]�������������̋�U��j�hx�h)d�    P���SVW���1E�3�P�E�d�    �e���P��!�E�}� t#�E�    �U��E�������   Ëe��E�����蠪���M�d�    Y_^[��]��������������������������������������������̋�U��E� ��M���U���E��]�����������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �}t�}u�T  �}t�}t�}t�}t
�}�F  j �	������E�    �}t�}u=�=� u4jh��	��"��u��   ��$"��������0�E�   �E�E̋M̃��M̃}���   �U���p�	�$�\�	� �Q��!�E�}t�UR��!� ��r��P��!�E�}t�MQ��!���L��R��!�E�}t�EP��!���%��Q��!�E�}t�UR��!���E������   �j �ͷ����Ã}� t��   ��   �}t�}t�}t��   �ğ���E؃}� u��   �E؁x\� uLhY  h(?j�pQ觞�����EȋU؋EȉB\�}� t�pQh� �U؋B\P輱������j�M؋Q\R�EP�5  ���E��}� u�L�M��Q�U�}t5�E��H;Mu*�U��E�B�M����M��tk��E�P\9U�r��ˋE��   �M�MċUă��Uă}�w�E�����	�$���	����x3�t	�E�   ��E�    �E��EЃ}� u!h�>j h�  hh>j�ͣ������u̃}� u.�����    j h�  hh>hT>h�>耻������������M�d�    Y_^[��]Ë���	D�	k�	�	��	 �I ˃	Ѓ	     ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    j 躣�����E�    �} u�E� ��E܋Q��!�E��E�   ��E���U܋P��!�E��E�   �}� t�}�t
�����M܉�E������   �j �2�����Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U�����	�$���	�E� ��MЋ�U�E؃��E��  �E���MЋ�U�E؃��E���   �E���MЋ�U�E؃��E���   �E���MЋ�U�E؃��E��   �����E��}� u�����  �M��Q\R�EP��  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h�>j h�  hh>j�џ������u̃}� u1脿���    j h�  hh>hd?h�>脷��������4  �E�P��!�E�}�u3��  �}� uj�����}� t
j �������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<�h�M��	�Uԃ��Uԡhl9E�}�M�k��U��B\�D    ���
�����MЉ�E������   ��}� t
j �K�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë��	��	T�	q�	7�	̇	 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��Q;Ut�E����E��tk�M9M�s�ًtk�U9U�s�E��H;Mu�E���3���]������������������������������������̋�U���P��!]�������������̋�U���'�����d]�����������������̋�U��������`]�����������������̋�U��E��]�����������������̋�U���$V��P��!�E�3Ƀ} ���M��}� uh�@j jDh@j��������u̃}� u0�ɻ���    j jDh@h@h�@�̳�����   �  �E�     �}� �_  h�� "�E�}� ut3�t	�E�   ��E�    �U��U�}� uh�?j jPh@j�{�������u̃}� u0�.����    j jPh@h@h�?�1������   ��   ht?�M�Q��!�E��}� ��   3�t	�E�   ��E�    �E܉E�}� uh�?j jVh@j��������u̃}� uD�$"P��������荺���0j jVh@h@h�?蔲�����$"P�������V�U�R��!�E�迢���E��E�Ph���";E�t
�M�Q��"j�UR�U���u�����    ����� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������̋�U��jj �EP�MQ��  ��]���������������������̋�U��jj �EPj ��  ��]�������̋�U��jj �EP�MQ�  ��]���������������������̋�U��jj �EPj �|  ��]�������̋�U��jj �EP�MQ�Z  ��]���������������������̋�U��jj �EPj �,  ��]�������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj ��  ��]��������������������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj �y  ��]��������������������̋�U��jh  �EP�MQ�G  ��]������������������̋�U��jh  �EPj �  ��]��������������������̋�U��jhW  �EP�MQ��  ��]������������������̋�U��jhW  �EPj �  ��]��������������������̋�U��jj�EP�MQ�  ��]���������������������̋�U��jj�EPj �\  ��]�������̋�U��jj �EP�MQ�:  ��]���������������������̋�U��jj �EPj �  ��]�������̋�U��jj �EP�MQ��   ��]���������������������̋�U��jj �EPj �   ��]�������̋�U����EP�M������M�芕���x t8�M��|����H�y�  u$jj �UR�EP�i   ���E�M�螶���E���E�    �M�芶���E��]��������������������������������̋�U��j �EP�p�����]�����������̋�U��j�h(�d�    P�����3�P�E�d�    �EP�M��2����E�    �M�M�M�譔���P�E�L#Mu;�} t�M�菔������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M�蓵���E��M�d�    Y��]��������������������������������������������������������������̋�U����} uh�Aj jdhXAj肔������u̋M�M��U�R�������E��E��H��   u$����� 	   �U��B�� �M��A����G  �-�U��B��@t"����� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6蛤���� 9E�t莤����@9E�u�M�Q�/�������u�U�R�p������E��H��  ��   �U��E��
+Hy!h�@j h�   hXAj��������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�)������E��q�}��t!�}��t�M����U������@�U���E�P��E��H�� t7jj j �U�R�<������E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P苑�����E�M�;M�t�U��B�� �M��A�����E%�   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M�蠞���E�    蛰���E�3Ƀ} �������������� u!h�Dj h  h�Dj衐������u̃����� uF�Q����    j h  h�DhdDh�D�Q�����ǅ ��������M������� �����  �E�������������Q��@��   ������P�Ԝ�����������������t-�������t$�������������������@������
ǅ���P�������H$�����х�uV�������t-�������t$�������������������@������
ǅ���P�������B$�� ���ȅ�tǅ ���    �
ǅ ���   �� ��������������� u!h0Cj h  h�Dj�,�������u̃����� uF�ܮ���    j h  h�DhdDh0C�ܦ����ǅ��������M��}���������U  3Ƀ} �������������� u!h�j h  h�Dj褎������u̃����� uF�T����    j h  h�DhdDh��T�����ǅ��������M�������������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���g  ������ �Z  �������� |%��������x���������A���������
ǅ����    ���������������������������B����������������������������  �������$�d�	�E�    �M�諌��P������R�1���������   ������P�MQ������R�t  ���E��������U���U����������؉�����u!hCj h�  h�Dj��������u̃����� uF蕬���    j h�  h�DhdDhC蕤����ǅ��������M��6���������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK����������	�$���	�E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP蝨�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�D������Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ��������Ĩ	�$���	�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ��������0�	�$���	�U���0  u�E�   �E��M���  tUǅ|���    �UR������f������������Ph   ������Q�U�R�l�������|�����|��� t�E�   �&�EP������f��x�����x����������E�   �������U��W  �EP��������t�����t��� t��t����y u�`��U��E�P�������E��P�M���   t&��t����B�E���t�����+����E��E�   ��E�    ��t����B�E���t�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������l����MQ�������E��U���  te�}� u�d��E��E�   �M���h�����l�����l�������l�����t��h������t��h�������h����ɋ�h���+M����M��[�}� u	�`��U��E���p�����l�����l�������l�����t��p������t��p�������p����ɋ�p���+E��E��  �MQ�9�������d����(�������   3�tǅ����   �
ǅ����    ��������`�����`��� u!h�Bj h�  h�Dj��������u̃�`��� uF蟦���    j h�  h�DhdDh�B蟞����ǅ��������M��@���������  ��  �U��� t��d���f������f����d�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  htBj�Ú�]  R������E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���X�����\����M��Ԅ��P�E�P�M�Q������R�E�P�M�Q��X���R��P��!�Ѓ��M���   t$�}� u�M�芄��P�U�R��P��!�Ѓ���������gu*�U���   u�M��U���P�E�P��Q��!�Ѓ��U����-u�M���   �M��U����U��E�P�������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�0�������H�����L����   �U���   t�EP��������H�����L����   �M��� tB�U���@t�EP轠��������H�����L�����MQ衠���������H�����L����=�U���@t�EP�{��������H�����L�����MQ�`�����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��M̋Ũ��U̅���@����D���t{�E��RP��D���Q��@���R�j�����0��T����E��RP��D���P��@���Q�|�����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �J  ���U�R������P�MQ�U�R�E�P�{  ���M���t$�U���u������P�MQ��<���Rj0��  ���}� ��   �}� ��   ǅ$���    �E���8����M܉�4�����4�����4�������4�������   ��8���f�f������������Pj��(���Q��0���R�}�������$�����8�������8�����$��� u	��0��� uǅ���������*�M�Q������R�EP��0���Q��(���R�z  ���V�����E�P������Q�UR�E�P�M�Q�T  �������� |$�U���t������P�MQ��<���Rj ��  ���}� tj�E�P�������E�    �v���������������M��#���������M�3��Ԣ����]�l�	h�	��	�	]�	i�	��	�	�	��	ߛ	ԛ	�	�	 �I �	̝	�	ם	�	 �w�	$�	d�	>�	Ξ	��	:�	�	��	�	7�	z�	.�	J�	%�	   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�}������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A�]��������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��E����U�
�E�f�A�]�������������������̋�S�܃������U�k�l$���   ���3ŉE��C��M��U��U�C��M��U����U��}�w@�E��$�@�	�E�   �4�E�   �+�E�   �"�E�   ��E�   ��K�   �E�    �}� ��   �U�P�K��Q�U�R�ӕ������ul�C�E�}�t�}�t�}�t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ�U�R�E�P��p���Q�����h��  �U�P�����ǅl���    �K�9t�=�� u�SR訓������l�����l��� u�C�Q�|�����M�3��������]��[��	#�	�	�	�	>�	5�	,�	���������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E�}� |,�}�~�}�t����M��U���y���E��o3�t	�E�   ��E�    �U��U��}� uh�Ej j9hHEj�t������u̃}� u+�<����    j j9hHEhEh�E�?����������E���]���������������������������������������������������̋�U��E��]�����������������̋�U���@���3ŉE��E�    �|���E��E�    �E�    �E�    �=� ��   hxF� "�Eԃ}� u3��  hhF�E�P��!�E��}� u3��  �M�Q��!��hTF�U�R��!P��!� �h<F�E�P��!P��!�$�hF�M�Q��!�E��U�R��!�,��=,� th F�E�P��!P��!�(��(�;M�th�,�;U�t]�(�P��!�EЋ,�Q��!�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W� �;M�t� �R��!�Eȃ}� t�UȉE�}� t*�$�;E�t �$�Q��!�Eă}� t
�U�R�UĉE��P��!�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��8�����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�Gj jhXGj� q������u̃}� u0賐���    j jhXGh@Gh�G趈�����   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E��M���Qh�   �U��R�=q����3��} ���E��}� uh�-j jhXGj�7p������u̃}� u0�����    j jhXGh@Gh�-�������   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E܋M���Qh�   �U��R�Dp������F��t3�t	�E�   ��E�    �U؉U�}� uh�Fj j hXGj�'o������u̃}� u0�ڎ���    j j hXGh@Gh�F�݆�����   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���MԋU���Rh�   �E��P�0o������-��t3�t	�E�   ��E�    �EЉE�}� uh<-j j*hXGj�n������u̃}� u-�ƍ��� "   j j*hXGh@Gh<-�Ʌ�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9<�s�<��U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�Fn����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�Gj jhXHj�l������u̃}� u0躋���    j jhXHh<Hh�G轃�����   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E�M���Qh�   �U��R�Hl����3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���M��U���Rh�   �E��P��k����3Ƀ} ���M��}� uh�-j jhXHj��j������u̃}� u0茊���    j jhXHh<Hh�-菂�����   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}�y����t&�M;Mrh�-j j+hXHj�+j������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E܋M���Qh�   �U��R�3j������-��t3�t	�E�   ��E�    �U؉U�}� uh<-j j>hXHj�i������u̃}� u-�Ɉ��� "   j j>hXHh<Hh<-�̀�����"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9<�s�<��M���U+U����E+EԋM���Qh�   �U+U��E�LPQ�Ii����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���E����E���t��E�+E������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�Gj jh .j��f������u̃}� u0胆���    j jh .h�Hh�G�~�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E�M���Qh�   �U��R�g����3��} ���E��}� uh�-j jh .j�f������u̃}� u0躅���    j jh .h�Hh�-�}�����   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���M��U���Rh�   �E��P�f������-��t3�t	�E�   ��E�    �E܉E�}� uh<-j jh .j��d������u̃}� u-蚄��� "   j jh .h�Hh<-�|�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9<�s�<��U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR�e����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�.j jhXHj�c������u̃}� u0�ʂ���    j jhXHh�Hh�.��z�����   �J  �} u\�U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U�E�Ph�   �M��Q�\c����3���  �} ��   �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U��E�Ph�   �M��Q��b����3҃} �U��}� uh�-j jhXHj��a������u̃}� u0裁���    j jhXHh�Hh�-�y�����   �#  �M�M��U�U��}�u5�E��M���E���U����U��E���E��t�M����M�t���y�)p����t&�U;Urh�-j j+hXHj�Da������u̋M��U���M���E����E��M���M��t�U����U�t�E���Et�} u�M�� �}� ��   �}�u�UU�B� �P   �?  �E�  �}�tI�}���t@�}v:�M��9<�s�<��U��	�E���E܋M�Qh�   �U��R�Wa������-��t3�t	�E�   ��E�    �U؉U�}� uh<-j j>hXHj�:`������u̃}� u-����� "   j j>hXHh�Hh<-��w�����"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9<�s�<��M���U+U����E+EԋM�Qh�   �U+U��E�LQ�o`����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��1l���MQ�UR�EP�MQ�M��]��P�.   ���E�M���~���E��]�������������������������̋�U����E�    �E��Q�U�j j �EP�MQ��"�E�}� u3���   �}� ~63�u2�����3��u��r#h��  �E�L Q�b����P�Iy�����E���E�    �U�U��}� u3��s�E�P�M�Q�UR�EP��"��u�H�F�} uj j j j j��M�Qj �U�R��!�E��!j j �EP�MQj��U�Rj �E�P��!�E��M�Q�.{�����E���]��������������������������������������������������������������������������̋�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�9{�����.�}���  t%3�u!h�Ij h�   hIj�L\������u̋�]��������������������������̋�U���$�} t�} v	�E�   ��E�    �E�E��}� uh�Gj jhJj��[������u̃}� u0�{���    j jhJh�Ih�G�s�����   �(  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9<�s�<��U��	�E+E��E�M���Qh�   �U��E�PQ�7Z����3���   3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E��M���Qh�   �U��R��Y������-��t3�t	�E�   ��E�    �U܉U�}� uh<-j jlhJj�X������u̃}� u-�mx��� "   j jlhJh�Ih<-�pp�����"   ��   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E�}� v�M����t�E���E�M���M��܋U����:u2�} t!�}s�  j�MQ�UR�EP�?s�����M���M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E؋M���Qh�   �U��R��V�����E�    �E�    �E�E��	�M���M�U����t4�M����/t�E����\u�U���U���E����.u�U�U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR�<r�����E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9<�s�<��M��	�U���UԋE���Ph�   �M��Q��U�����}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR�q�����}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R�[q�����   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR� q�����}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9<�s
�<��E��	�M(���MЋU���Rh�   �E$��P��T����3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9<�s�<��M��	�U���ŰE���Ph�   �M��Q�kT�����} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���EȋM���Qh�   �U��R�T�����} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9<�s
�<��E��	�M ���MċU���Rh�   �E��P�S�����}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9<�s�<��M��	�U(���U��E���Ph�   �M$��Q�=S����3҃} �U��}� u!hxKj h�   h�Jj�4R������u̃}� u3��q���    j h�   h�Jh�JhxK��i�����   �   �}� tw3�t	�E�   ��E�    �U��U܃}� u!h�Jj h�   h�Jj�Q������u̃}� u0�gq���    j h�   h�Jh�Jh�J�gi�����   ��7q��� "   �"   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���]��������̋�U����} |�}}	�E�   ��E�    �E��E��}� u"hXMj jqh�Lj�O������u�uH���}� u.�/o���    j jqh�Lh�LhXM�2g��������   �}�t�U���t	�E�    ��E�   �E�E�}� u"h�Kj jvh�Lj� O������u��G���}� u+�n���    j jvh�Lh�Lh�K�f��������/�}�u�U��p���E��p��M��U�E��p��E���]������������������������������������������������������������������������������������������̋�U����} |�}}	�E�   ��E�    �E�E��}� u%hXMj h�   h�Lj��M������u��F���}� u0�m���    j h�   h�Lh�MhXM�e����������c�}�u�U��|��Q�E��|��M��}�uj��@"�U��|��'�}�uj��@"�M��|���U�E��|��E���]��������������������������������������������������������������̋�U��Q���E��M���E���]������������������̋�U���]����̋�U��j�h(�h)d�    P���PP  �3K�����1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�4M����ƅ���� h�  j ������Q�M����3�f������h�  j ������P��L����ƅЯ�� h�  j ��ѯ��Q��L�����} |�}|����*  �E�    �}��   hl��"����   j h  h�Lh Th�Sj
h   ��п��R�EP�<e����P�aZ����h�S��"�} t�M�������
ǅ����|S������R��"hpS��"��п��P��"h����"�2D��ǅ���������=  �} ��   ǅ̯��    ��j�����ȯ����j���     �UR�EPh�  h   ��Я��Q�Bg������̯����̯�� }*j h*  h�Lh Th��j"j�mj���R�E���� �]j����ȯ�����̯�� }8j h-  h�Lh Th�Rh�h   ��Я��R�tk����P�#Y�����}uV�} tǅ�����R�
ǅ�����Rj h2  h�Lh Th�Q������Ph   ��п��Q�k����P��X����j h4  h�Lh ThHQ��Я��Rh   ��п��P�%B����P�X�����}u�M��p���t8j h9  h�Lh Th�Ph�Ph   ��п��P��A����P�@X����j h:  h�Lh Th�Ph��h   ��п��Q�A����P�X�����} ��   ǅį��    ��h�����������h���     ��п��P�MQ�URh|Ph�  h   ������P�oL������į����į�� }*j hA  h�Lh Th��j"j�rh���Q�C���� �bh�����������į�� }8j hD  h�Lh Th�h�h   ������P�yi����P�(W�����:j hH  h�Lh ThP��п��Qh   ������R�=i����P��V����ǅ����    ǅ����    j�������Ph   ������Q������R�\����������j hM  h�Lh ThhOj"j������P��B���� ������ t8j hO  h�Lh Th�Nh�Mh   ������Q�Jh����P�DV�����=� u�=� �#  ǅ����    ǅ����    j��H�����E�   ����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j��X����Ã����� �D  �=� t?ǅ����    ������R������P�MQ������tǅ����   ������������������ ��   �E��p���t>�U�<�|��t1j ������P������Q��I����P������R�E��|�Q��"�U��p���t������Q��"�U��p���twƅп�� �} t9j h�  h�Lh Th�Sj
h   ��п��Q�UR��^����P��S������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�=h�����������E������   ��}uhl��("Ë������M�d�    Y_^[�M�3��h����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hX�h)d�    P���\�  �A�����1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q�C����3�f������h�  j ������P��B����ƅ���� h�  j ������Q��B����3�f��Џ��h�  j ��ҏ��P�B�����} |�}|����.  �E�    �}��   hl��"����   j h�  h�Lhh[h[j
h   ��Я��Q�UR�T����P�-P����h�Z��"�} t�E������
ǅ����Z�����Q��"hlZ��"��Я��R��"hhZ��"��9��ǅ���������A  �} ��   �`��� ��ȏ���`���     �MQ�URh�  h   ��Џ��P�^X������̏����̏�� }*j h  h�Lhh[h��j"j�C`���Q�;���� �3`����ȏ�����̏�� }8j h  h�Lhh[h�Yh�h   ��Џ��P��`����P��N�����}uV�} tǅ���|Y�
ǅ���PYj h  h�Lhh[h�X�����Qh   ��Я��R�`����P�N����j h  h�Lhh[hX��Џ��Ph   ��Я��Q� 8����P�cN�����}u�U��p���t8j h  h�Lhh[h�Wh�Wh   ��Я��Q�7����P�N����j h  h�Lhh[hXWhhZh   ��Я��R�{7����P��M�����} ��   ǅď��    �^��� �������^���     ��Я��Q�UR�EPh<Wh   h   ������Q�);������ď����ď�� }*j h  h�Lhh[h��j"j�H^���R�9���� �8^�����������ď�� }8j h  h�Lhh[h�h�h   ������R�_����P��L�����:j h"  h�Lhh[h�V��Я��Ph   ������Q��^����P��L����ǅ����    j h(  h�Lhh[h Vj"jj�������Rh   ������Pj �*`����P�8���� ������������ t8j h*  h�Lhh[h8Uh�Th   ������Q�^����P�/L�����=� u�=� �#  ǅ����    ǅ����    j��>�����E�   ����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j��N����Ã����� �g  �=� t?ǅ����    ������R������P�MQ������t������������ǅ����   ������ �  �E��p����[  �U�<�|���J  �E��|�Q�H"����������t�Jj ������R������P�-?����P������Q�U��|�P��"��t��   �$"��t��   ǅ���    j h{  h�Lhh[hHTj"jj�������Qh   �����R�����P�g]����P��5���� ���������� t>�����Pt5j ������Q������R�z>������P������P�M��|�R��"�@����� v������������j ������Q�����R�����P�M��|�R��"�E��p���t������R��"�E��p���ty3�f��Я���} t9j h�  h�Lhh[h[j
h   ��Я��P�MQ�&M����P�H������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ�]�����������E������   ��}uhl��("Ë������M�d�    Y_^[�M�3���\����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���@���3ŉE��E�    �0?���E��E�    �E�    �E�    �=4� ��   hxF� "�Eԃ}� u3��  h�[�E�P��!�E��}� u3��  �M�Q��!�4�hTF�U�R��!P��!�8�h<F�E�P��!P��!�<�h�[�M�Q��!�E��U�R��!�D��=D� th F�E�P��!P��!�@��@�;M�th�D�;U�t]�@�P��!�EЋD�Q��!�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�8�;M�t�8�R��!�Eȃ}� t�UȉE�}� t*�<�;E�t �<�Q��!�Eă}� t
�U�R�UĉE�4�P��!�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��XX����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} u3��k  3��} ���E��}� uh�\j j7h(\j�)4������u̃}� u0��S���    j j7h(\h\h�\��K�����   �  �} t�U;U��   �EPj �MQ�4����3҃} �U��}� uh�[j j=h(\j�3������u̃}� u-�RS���    j j=h(\h\h�[�UK�����   �~�M;M҃��U�uh�[j j>h(\j�>3������u̃}� u-��R��� "   j j>h(\h\h�[��J�����"   ��   ��MQ�UR�EP�@����3���]�������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����������������������̋�U���D�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� u!h�j h�   h�\j��1������u̃}� u1�Q���    j h�   h�\h�\h��I��������Z  3Ƀ} ���M̃}� u!h�<j h�   h�\j�u1������u̃}� u1�(Q���    j h�   h�\h�\h�<�(I���������   �E�E��M��AB   �U�E�B�M�U��E��@����M�Qj �UR�E�P��Q�����E��} u�E��   �M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj ��H�����EċE�H���M��U�E��B�}� |!�M�� 3�%�   �E��M����E���M�Qj �H�����E��E���]��������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�E������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�:������]����������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�6>������]������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�<������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�S9������]��������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�t=������]����������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��;������]��������������������̋�U��Q�E�E��M�Q�UR�36������]����������������̋�U��Q�E�E��M�Q�UR�0������]����������������̋�U��Q�E�E��M�Q�UR�EP�\0������]������������̋�U��Q�E�E��M�Q�UR�EP�&E������]������������̋�U��Q�} t��}��E�P�V  ���M��} t
��  �U���]��������������������������̋�U�����}��E�P�
  ���E��=` t�]�M�Q��  ��E���E���]�������������������������������̋�U��QV�}���=` t�E�P�  �����w  ����M�Q�  ��^��]�������������������������������̋�U����} t^��}��E�P��  ���E�M#M�U��#U�ʉM��E�;E�t'�M�Q�Z  ��f�E��m���}��U�R�  ���E��E�M���} t)�=` t�UR�EP��  ���M��	�U�    �   ��]��������������������������������������������̋�U��E%����P�MQ�*����]��������������������̋�U�����}��E�P��  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�`  ��f�E��m���}��U�R�  ���E�=` tB�EP�MQ��  ���E�U�#P]�E�#P];�t�E�E�   ����E�E����E��]������������������������������������������������̋�U����} 	 u>�}�u8��}��E�%=  ==  u$�=` t�]��M�����  ���  u�;��7j h[  h ^h�]hX]�U������R�EPj �@����P�8������]��������������������������������������̋�U����S,��� �E�����!���R	  �}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]�������������������������̋�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]��������������������������������������������������������������������������������������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��������������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�������������������������������������̋�U��Q�Y&���E��E�P�)  ����]������������������̋�U��Q�]��e���U��E�P��  ����]��������������̋�U����E%�E�]��M�Q�   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R��  ���E��E�P��"�����]��M�Q�2   ����]�������������������������������������������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]��������������������������������������������������������������������������������������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]��������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]��������������������������������������������̋�U��Q�E��  �E�P�������]�������������������̋�U���]����̋�U���]����̋�U����D+���E��E��Hp����Ƀ��M��U�U��E����E��}�wC�M��$��
�U��Bp���M��Ap�   �U��Bp����M��Ap�   �   �H������u3�t	�E�   ��E�    �E�E�}� u!h�`j h�   h`j�"������u̃}� u.��>���    j h�   h`h�_h�`��6���������E���]Ðo
j
B
V
�����������������������������������������������������������������������̋�U��j�h��h)d�    P��SVW���1E�3�P�E�d�    �=� �tAj�������E�    h �h��y:�������E������   �j�0����ËM�d�    Y_^[��]�����������������������������������������������̋�U��j�h��h)d�    P��SVW���1E�3�P�E�d�    �} ��   j�0�����E�    �E�x t.�M�QR�("��u�E�x �tj�M�QR�0�����E������   �j��/����ËE�8 tcj�������E�   �M�R��7�����E�8 t#�M��: u�E�8 �t�M�R�}A�����E������   �j�^/����ËE� 𭺋M�A�j�UR��/�����M�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��EP�z����]�������������̋�U����E�    �} |�}�} u3��  he  h�`jjj�:�����E��}� u�;���    3��  hj  h�`jjh�   �o:�����M���U��: u j�E�P��.�����F;���    3��8  hp  h�`jjh   �':�����E��M��U��Q�}� u0j�E��Q�.����j�U�R�.������:���    3���   h ��E��Q�P  ���UR�EP�M��R�z  ����u3�E��Q�5�����U��P�s?����j�M�Q�!.�����E�    �x�U��BP�M���BP��������tDj�M��QR��-�����E��Q�I5�����U��P�?����j�M�Q��-�����E�    ��U��B�    �M��Q�   �E���]���������������������������������������������������������������������������������������������������������������������������������̋�U��VW�} t0�} t*�E;Et"�u�6   �}�M�    �UR�M3����_^]�������������������������������̋�U��EP�MQ�(����]���������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�    �s$���E�h�  h�`jjj�7�����E�}� u�8���    3��   �%-���0���E�M��Ql��E�M��Qh�Pj�G�����E�    �E�Q�V2�����E������   �j�	+�����j������E�   �U�BP�"�E������   �j��*����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������̋�U���T/��]����̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �EԉE؃}� u!hHaj h&  h`j�E������u̃}� u0��6���    j h&  h`h0ahHa��.����3��  �}"���E��b+���U܋Bp���M܉Ap�E�    h1  h�`jjh�   �5�����E�}� �  j�b�����E�   �U܋BlP�M�Q��������E�    �   �j�)����Ã}� ��   �UR�EP�M�Q��  ���E��}� ��   �} thL��UR��������t
�L�   j�������E�   �E�P�M܃�lQ�_2�����U�R��0�����E܋Hp��u$�H���u�E܋HlQh��)2�����
  �E�    �   �j�W(�������U�R�w0�����E�P�C:�����E������   ��M܋Qp���E܉PpËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U������   ��������   �������   �h�]���������������������̋�U���   ���3ŉE��} tC�} t�EP�MQ�UR�  ����T�����E���M�TH��T�����T����E��|  ǅd���   ǅh���    �} �O  �M���L�'  �E�H��C�  �U�B��_�  �M��`���h|b��`���R�X������\�����\��� t"��\���+�`�����X���t��\������;u3���  ǅl���   ���l�������l�����l���N��X���Q��`���R��l���k����^Q�)������u"��l���k����^P�O����9�X���u�뚋�\�������\���hxb��\���R�"������X�����X��� u��\������;t3��$  ��l���|j h�  h`hLbh�a��X���R��\���Ph�   ��p���Q�h����P�H!������X���Ƅp��� ��p���P��l���Q�UR��  ����t��h�������h�����\����X�����`�����`������t��`�������`�����`�������7�����h��� t�MQ��  ����P����
ǅP���    ��P����U��  �EPj j h�   ��p���Q�UR��,�����E��}� ��   ǅl���    ���l�������l�����l���|��l��� tn��l������U�D
HP��p���Q��������t;��p���R��l���P�MQ�  ����t��h�������h����
ǅd���    ���h�������h����l�����d��� t�MQ��  ���E��0��h��� t�UR�  ����L����
ǅL���    ��L����E���MQ�  ���E��E��M�3���3����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ���3ŉE�ǅX���    ǅT���    ������D�����D����  ��l���ǅH���   �MQ��@���R��L���Ph�   ��p���Q�UR�g*������u3��  �E���M�THR��p���P�j������u�M���U�D
H�a  ��p���P����������T���h�  h�`j��T���Q�w������X�����X��� u3��  �U���E�LH��8����U�E�L���<���j�Uk��E�L$Q��0���R�a�����E�H��\���j h  h`hch�b��p���R��T�����P��X�����Q�/����P��������X������E���M�TH��L����E�M�T�j��L���R�Ek��M�T$R�������}�
  �E��@����H��H�����l����L���T����(�����,���ǅ`���    ���`�������`�����`���;�H�����   �U��`�����l����R;�uJ��`��� t=��`�����l������D���l�����A��`�����l�����(����Ћ�,����L��]�V��`�����l����ЋT���d�����h�����`�����l�����(�������,����T���d�����(�����h�����,����#�����`���;�H�����   j�E�HQ�U�BP��8���Qjh@_jj �K���� ����   ǅ$���    ���$�������$�����$���s$��$�����E8������  ��$���f��U8�����h�   ���P��8���Q�������u��l����B   ���l����@    ���l����A    ��l����E�H�
�U��l����H���   �}u�U��@����B�MQ�Uk����^�Ѓ���tG�M���U��8����D
Hj��X���Q������U�E��<����L��U��\����B3��   ��8���L�t{�M���U�D
PP�("��uc3�uj j h[  h`j��
������u�j�E���M�TPR�.����j�E���M�TTR������E���M�DL    ��X��� t��X����   �E���M��X����TP�E���M�DH�M�3���-����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�    �E�    �E�    �E�U  ht  h�`j�E�P������E�}� u3��  �M���M��U���U��E��  �M��   �E�   �	�U����U��E����M�THRh�4�E�k����^Qj�U�R�E�P�)�����}�}kj h�  h`hpch4chxb�M�Q�U�R� ����P�������E������M�THR�E����M�THR�{������t�E�    �  �}� ��   �E�xP tD�M�QPR�("��u33�uj j h�  h`j�������u�j�U�BPP�������M�yT tD�U�BTP�("��u33�uj j h�  h`j�[������u�j�E�HTQ������U�BT    �E�@L    �M�U�QP�E�M��HH�E���   ��   j�U�R�c�����E�xP tD�M�QPR�("��u33�uj j h�  h`j��������u�j�U�BPP������M�yT tD�U�BTP�("��u33�uj j h�  h`j�������u�j�E�HTQ�������U�BT    �E�@L    �M�AP    �U�BH    �E�@h�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����   ���3ŉE������   �E�E��(�E��M�� �M�U��,�U��E�   �E��   �E��E��   �E�    �} u3��-  �} t�} u3��  �M���Cuv�E�H��ukj h�  h`h�dh�dh�d�UR�EP��%����P�t�����} t3ɋUf�
3��Mf�A3ҋEf�P�} t	�M�    �E�  �UR������E��}��   s0�EP�M�Q���������  �UR�E�P���������   ǅ@���    ǅD���    �MQ��H���R�������t3��  ��H���P�M�Q��H���R�������u3���   �E��H�U��
��H���P�M�Q�U�R�k	�����E���t�}��   s�U��@����E���D����
ǅ@���+�j h�  h`h�dh d��D�����Q��@���R�E�P�M�Q�* ����P�
�����} tj�U�R�EP�:�����} tj�M�Q�UR�"����j h  h`h�dh�c�E�P�MQ�UR��#����P������E��M�3��#&����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�]�������̋�U����E�E��E�    �	�M����M��U�;U}A�E����E�j h  h`h�fhe�M��Q�R�EP�MQ������P�t������E�    ��]��������������������������������������������̋�U���h�   j �EP�)�����M���u3���  �E���.uX�U�B��tMj h*  h`h�jh�ij�M��Qj�U�   R�������P������Eƀ�    3��e  �E�    �	�M����M�h�i�UR��������E��}� u����1  �EE���M��}� uI�}�@sC�U���.t:j h8  h`h�jh�h�E�P�MQj@�UR�C�����P�#�����   �}�uI�}�@sC�E���_t:j h;  h`h�jh�g�M�Q�URj@�E��@P�������P�������_�}�uT�}�sN�M���t	�U���,u=j h>  h`h�jh�f�E�P�MQj�U�   R������P�w���������)�E���,u��M���u��U��E�L�M����3���]����������������������������������������������������������������������������������������������������������������������������������������̋�U��j hT  h`hxkh�j�EP�MQ�UR������P������E�H@��t�U��@Rh�jj�EP�MQ�W������U���   ��t!�M���   Qh�jj�UR�EP�(�����]����������������������������������������������̋�U����EP�M������M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M��:���P�.   ��$�E�M��s���E��]�������������������������̋�U��� �} ~,�EP�MQ�%  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R��!�E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R�:����P�~�����E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R��!��u
�Y  �T  j j �E�P�M�Q�UR�EP��"�E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR��"��u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�3 ����P�w�����E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ��"��u�V�T�}  u+j j j j �U�R�E�Pj �M$Q��!�E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P��!�E��}� t�M�Q�@�����U�R�4�����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U����EP�M������M��J�����U���   �P�� �  �M�M��v���E��]����������������������������̋�U��j �EP������]�����������̋�U��h  �EP�����]�������̋�U��h  �EP������]�������̋�U��j�EP������]����������̋�U��j�EP�����]����������̋�U��j�EP�����]����������̋�U��j�EP�v����]����������̋�U��j�EP�V����]����������̋�U��j�EP�6����]����������̋�U��h�   �EP�����]�������̋�U��h�   �EP������]�������̋�U��j�EP������]����������̋�U��j�EP�����]����������̋�U��j�EP�����]����������̋�U��j�EP�v����]����������̋�U��h  �EP�S����]�������̋�U��h  �EP�3����]�������̋�U��hW  �EP�����]�������̋�U��hW  �EP������]�������̋�U��h  �EP������]�������̋�U��h  �EP�����]�������̋�U��j �EP�����]����������̋�U��j �EP�v����]����������̋�U���E=�   ���]������������̋�U��Qh  �EP�2������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�B������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ����������������������������XY�$�����������XY�$�����������XY�$����������̋�U���SVWd�5    �u��E�3
j �EP�M�Q�UR� ���E�H����U�Jd�=    �]��;d�    _^[��]� ����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�^���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ����� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ����� �E�_^[�E���]��������������������̋�U��E�HQ�U�B(Pj �M�QR�\�����]� �����������������������̋�U����E�    �E�5
����M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ�
����E�E�d�    �E��]����������������������������������̋�U��Q��E�H3M���j �MQ�U�BP�M�QRj �EP�M�QR�EP����� �E��E���]��������������������̋�U���8S�}#  u�.6
�M��   ��   �E�    �Eܠ6
����M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M��C������   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]��������������������������������������������������������������������̋�U��QS��E�H3M�~���M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ��	���� �U�z$ u�EP�MQ��	��j j j j j �U�Rh#  �,������E��]�c�k ��   [��]���������������������������������������������������̋�U��Q�} �E�HSV�pW�M�����|8����u�����E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v������M�_��^��[��]��������������������������������̋�U��EV�u��������   �N�������   ��^]��������������������̋�U����������   ��t�M9t�@��u��   ]�3�]�������������������̋�U��V�����u;��   u�����N���   ^]��������   �x t�H;�t���x u�^]������V�P^]�������������������������̋�U����EP�M��q����M$Q�U R�EP�MQ�UR�EP�MQ�M������P�2   �� �E�M�����E��]�����������������������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP��!�E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP� �����P�d	�����E���E�    �M�M��}� u3��a�U���Rj �E�P�|������M�Q�U�R�EP�MQj�UR��!�E��}� t�EP�M�Q�U�R�EP��"�E��M�Q�[�����E���]�����������������������������������������������������������������������̋�U��Q�E�x  toj?hdljhd  j������E��}� u
�   �   �MQ�U�R��   ����t!�E�P�!����j�M�Q�  �����   �}�U�ǂ�      ��E�P��E���   P�tJ�M���   �´   R�("��u0�E���   ���    hlj jOh�kj�0�������u̋E�M����   3���]����������������������������������������������������������������̋�U����E�    �E�HB�M��U�BD�E��} u�����  �M�M��E�    �U��Rj1�E�Pj�M�Q�������E�E�U��Rj2�E�Pj�M�Q������E�E�U��Rj3�E�Pj�M�Q������E�E�U��Rj4�E�Pj�M�Q�q�����E�E�U��Rj5�E�Pj�M�Q�P�����E�E�U��Rj6�E�Pj�M�Q�/�����E�E�URj7�E�Pj�M�Q������E�E�U�� Rj*�E�Pj�M�Q�������E�E�U��$Rj+�E�Pj�M�Q�������E�E�U��(Rj,�E�Pj�M�Q������E�E�U��,Rj-�E�Pj�M�Q������E�E�U��0Rj.�E�Pj�M�Q�l�����E�E�U��4Rj/�E�Pj�M�Q�K�����E�E�U��Rj0�E�Pj�M�Q�*�����E�E�U��8RjD�E�Pj�M�Q�	�����E�E�U��<RjE�E�Pj�M�Q�������E�E�U��@RjF�E�Pj�M�Q�������E�E�U��DRjG�E�Pj�M�Q������E�E�U��HRjH�E�Pj�M�Q������E�E�U��LRjI�E�Pj�M�Q�d�����E�E�U��PRjJ�E�Pj�M�Q�C�����E�E�U��TRjK�E�Pj�M�Q�"�����E�E�U��XRjL�E�Pj�M�Q������E�E�U��\RjM�E�Pj�M�Q�������E�E�U��`RjN�E�Pj�M�Q������E�E�U��dRjO�E�Pj�M�Q������E�E�U��hRj8�E�Pj�M�Q�}�����E�E�U��lRj9�E�Pj�M�Q�\�����E�E�U��pRj:�E�Pj�M�Q�;�����E�E�U��tRj;�E�Pj�M�Q������E�E�U��xRj<�E�Pj�M�Q�������E�E�U��|Rj=�E�Pj�M�Q�������E�E�U�   Rj>�E�Pj�M�Q������E�E�U�   Rj?�E�Pj�M�Q������E�E�U�   Rj@�E�Pj�M�Q�l�����E�E�U�   RjA�E�Pj�M�Q�H�����E�E�U�   RjB�E�Pj�M�Q�$�����E�E�U�   RjC�E�Pj�M�Q� �����E�E�U�   Rj(�E�Pj�M�Q�������E�E�U�   Rj)�E�Pj�M�Q������E�E�U�    Rj�E�Pj�M�Q������E�E�U�¤   Rj �E�Pj�M�Q�p�����E�E�U�¨   Rh  �E�Pj�M�Q�I�����E�E�U�°   Rh	  �E�Pj �M�Q�"�����E�E�U�E����   �M���   Qj1�U�Rj�E�P�������E�E�M���   Qj2�U�Rj�E�P�������E�E�M���   Qj3�U�Rj�E�P������E�E�M���   Qj4�U�Rj�E�P������E�E�M���   Qj5�U�Rj�E�P�b�����E�E�M���   Qj6�U�Rj�E�P�>�����E�E�M���   Qj7�U�Rj�E�P������E�E�M���   Qj*�U�Rj�E�P�������E�E�M���   Qj+�U�Rj�E�P�������E�E�M���   Qj,�U�Rj�E�P������E�E�M���   Qj-�U�Rj�E�P������E�E�M���   Qj.�U�Rj�E�P�f�����E�E�M���   Qj/�U�Rj�E�P�B�����E�E�M���   Qj0�U�Rj�E�P������E�E�M���   QjD�U�Rj�E�P�������E�E�M���   QjE�U�Rj�E�P�������E�E�M���   QjF�U�Rj�E�P������E�E�M���   QjG�U�Rj�E�P������E�E�M��   QjH�U�Rj�E�P�j�����E�E�M��  QjI�U�Rj�E�P�F�����E�E�M��  QjJ�U�Rj�E�P�"�����E�E�M��  QjK�U�Rj�E�P�������E�E�M��  QjL�U�Rj�E�P�������E�E�M��  QjM�U�Rj�E�P������E�E�M��  QjN�U�Rj�E�P������E�E�M��  QjO�U�Rj�E�P�n�����E�E�M��   Qj8�U�Rj�E�P�J�����E�E�M��$  Qj9�U�Rj�E�P�&�����E�E�M��(  Qj:�U�Rj�E�P������E�E�M��,  Qj;�U�Rj�E�P�������E�E�M��0  Qj<�U�Rj�E�P������E�E�M��4  Qj=�U�Rj�E�P������E�E�M��8  Qj>�U�Rj�E�P�r�����E�E�M��<  Qj?�U�Rj�E�P�N�����E�E�M��@  Qj@�U�Rj�E�P�*�����E�E�M��D  QjA�U�Rj�E�P������E�E�M��H  QjB�U�Rj�E�P�������E�E�M��L  QjC�U�Rj�E�P������E�E�M��P  Qj(�U�Rj�E�P������E�E�M��T  Qj)�U�Rj�E�P�v�����E�E�M��X  Qj�U�Rj�E�P�R�����E�E�M��\  Qj �U�Rj�E�P�.�����E�E�M��`  Qh  �U�Rj�E�P������E�E�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u�W  j�E�HQ�������j�U�BP�������j�M�QR������j�E�HQ������j�U�BP������j�M�QR������j�E�Q�r�����j�U�B P�a�����j�M�Q$R�P�����j�E�H(Q�?�����j�U�B,P�.�����j�M�Q0R������j�E�H4Q������j�U�BP�������j�M�Q8R�������j�E�H<Q�������j�U�B@P�������j�M�QDR������j�E�HHQ������j�U�BLP������j�M�QPR������j�E�HTQ�s�����j�U�BXP�b�����j�M�Q\R�Q�����j�E�H`Q�@�����j�U�BdP�/�����j�M�QhR������j�E�HlQ������j�U�BpP�������j�M�QtR�������j�E�HxQ�������j�U�B|P�������j�M���   R������j�E���   Q������j�U���   P������j�M���   R�y�����j�E���   Q�e�����j�U���   P�Q�����j�M���   R�=�����j�E���   Q�)�����j�U���   P������j�M���   R������j�E���   Q�������j�U���   P�������j�M���   R�������j�E���   Q������j�U���   P������j�M���   R������j�E���   Q�u�����j�U���   P�a�����j�M���   R�M�����j�E���   Q�9�����j�U���   P�%�����j�M���   R������j�E���   Q�������j�U���   P�������j�M���   R�������j�E���   Q�������j�U���   P������j�M���   R������j�E���   Q������j�U��   P�q�����j�M��  R�]�����j�E��  Q�I�����j�U��  P�5�����j�M��  R�!�����j�E��  Q������j�U��  P�������j�M��  R�������j�E��   Q�������j�U��$  P������j�M��(  R������j�E��,  Q������j�U��0  P������j�M��4  R�m�����j�E��8  Q�Y�����j�U��<  P�E�����j�M��@  R�1�����j�E��D  Q������j�U��H  P�	�����j�M��L  R�������j�E��P  Q�������j�U��T  P�������j�M��X  R������j�E��\  Q������j�U��`  P������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �E�    �E�E��E�    �M�y u�U�z �  jeh`mjjPj�������E�}� u
�   ��  �E���   �   �}��jqh`mjj��������E�}� uj�M�Q�H������   �z  �U��    �E�x �:  j}h`mjj�������E��}� u&j�M�Q�������j�U�R��������   �"  �E��     �M�Q>�U��E�Pj�M�Qj�U�R������E�E�E��Pj�M�Qj�U�R������E�E�E��Pj�M�Qj�U�R�n�����E�E�E��0Pj�M�Qj�U�R�M�����E�E�E��4Pj�M�Qj�U�R�,�����E�E�t0�E�P������j�M�Q������j�U�R����������;  �E�HQ�  ���@�E�    �U䡠���M����Q�E����H�U����B0�M����Q4�E��    �}� t	�M��   ��E�    �E�    �E���U���    tA�E���   Q�("��u-�U���    w!hmj h�   h�lj���������u̋M���    t<�U���   P�("��u(j�M���   R�������j�E���   Q��������U�E����   �M�U쉑�   �E�M䉈�   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�   �E�;��tj�U�P�������M�Q;��tj�E�HQ��������U�B;��tj�M�QR��������E�H0;��tj�U�B0P�������M�Q4;��tj�E�H4Q������]�����������������������������������������������������̋�U���VW�E�    �E�E��E�    �M�y u�U�z �W  jSh`njjPj�������E�}� u
�   ��  jYh`njj�r������E��}� uj�E�P��������   ��  �M��    �U�z �d  jeh`njj�(������E�}� u&j�E�P������j�M�Q�������   �s  �U��    �E�H8�M��E�    �U��Rj�E�Pj�M�Q�@�����E�E�U��Rj�E�Pj�M�Q������E�E�U��Rj�E�Pj�M�Q�������E�E�U��Rj�E�Pj�M�Q�������E�E�U��Rj�E�Pj�M�Q������E�E�U�� RjP�E�Pj�M�Q������E�E�U��$RjQ�E�Pj�M�Q�z�����E�E�U��(Rj�E�Pj �M�Q�Y�����E�E�U��)Rj�E�Pj �M�Q�8�����E�E�U��*RjT�E�Pj �M�Q������E�E�U��+RjU�E�Pj �M�Q�������E�E�U��,RjV�E�Pj �M�Q�������E�E�U��-RjW�E�Pj �M�Q������E�E�U��.RjR�E�Pj �M�Q������E�E�U��/RjS�E�Pj �M�Q�r�����E�E�U��8Rj�E�Pj�M�Q�Q�����E�E�U��<Rj�E�Pj�M�Q�0�����E�E�U��@Rj�E�Pj�M�Q������E�E�U��DRj�E�Pj�M�Q�������E�E�U��HRjP�E�Pj�M�Q�������E�E�U��LRjQ�E�Pj�M�Q������E�E�t@�U�R�a�����j�E�P������j�M�Q������j�U�R�y������   �b  �E�HQ�  ����   ����}��U���   �M���E���   �U�A�B�M���   �E�J�H�U���   �M�P0�Q0�E���   �U�A4�B4�M��   �}� t	�U��   ��E�    �E�    �E���E���    tA�M���   R�("��u-�E���    w!hnj h�   h�mj�!�������u̋U���    t<�E���   Q�("��u(j�U���   P�G�����j�M���   R�3������E�M䉈�   �U�E����   �M�U艑�   3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�  �E�H;��tj�U�BP��������M�Q;��tj�E�HQ�������U�B;��tj�M�QR�������E�H;��tj�U�BP�|������M�Q;��tj�E�HQ�]������U�B ;��tj�M�Q R�>������E�H$;��tj�U�B$P�������M�Q8;��tj�E�H8Q� ������U�B<;��tj�M�Q<R��������E�H@;��tj�U�B@P��������M�QD;��tj�E�HDQ�������U�BH;��tj�M�QHR�������E�HL;��tj�U�BLP�e�����]�����������������������������������������������������������������������������������������������������������̋�U��������E��E��Hl�M��U�;�t�E��Hp#H�u������E������]�����������������������������̋�U���]����̋�U��������E��E��Hl�M��U�;�t�E��Hp#H�u�W����E��U����   ��]�������������������������̋�U��h��EP�MQ������]��������������������̋�U���<���3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q���������t	�E�    ��U�R��������E�   �Z  �E�P�M�Q�,������U�U؋E�HQ�U�R�C�������t	�E���E�M�U�A+B9E�}�M�Q�������E�    �E�   ��   �U�E�;Bk�M�Q�U�R軻�����E؉E�M�Q+U�UċE�P�M�Q�������U�BP�M�Q�������U�B��P�M�Q��������E�    �E�   �~�U�E�;|B�M�Q��������U܁�   ��U܋E�HQ�U�R�������E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�g������E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3�������]������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ��������u�U�R�EP�������E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������������������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]��������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P��������E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�������E��ȋE���]������������������������������������������������������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]����������������̋�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]����������������������������������̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�����������������������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]������������������������������������������������������������������̋�U��h,��EP�MQ�L�����]��������������������̋�U������3ŉE��E�    �E�H
���  f�M��U�B
% �  f�E�M�Q�U�E�H�M�U����E�j@�M�Q�L�������t�E�   �f�U�f��f�U��E�=�  u�E�   �M�U�Q�E�M��U��E�ЋMf�Q�E��M�3��������]��������������������������������������������������������������̋�U���   ���3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!hyj h�   hhxj譺������u̃}� u0�`����    j h�   hhxhDxhy�`�����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$�4v
�U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p�����tv
�$�dv
�E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h������v
�$��v
�E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�����w
�$��v
�E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�������}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�K�����f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3�������]Ë��m
�n
Uo
�o
�p
�q
�q
�r
fr
s
$t
�s
.o
o
%o
@o
  ��p
}p
�p
  �{q
rq
�q
  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U������3ŉE������`�E��} u�   �} }�M�ىM�0���`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP�������눋M�3��s�����]�����������������������������������������������������������̋�U���L���3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q������f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R�٨����f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3��B�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]������������������������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]���������������������������̋�U������3ŉE��EPj j j �MQ�UR�EP�M�Q������ �E�UR�E�P�������E��}�u	�M���M�E�M�3��������]��������������������������������������̋�U���x���3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h�zh�zhXzhLzj�U��R�������P譳�����E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h�zh�zh�yh�yj�U��R������P�N������E�@�E�    �   �}�   �uK�}� uEj h�   h�zh�zh�yh�yj�M��Q�H�����P��������U�B�E�    �Cj h�   h�zh�zh8yh0yj�E��P������P貲�����M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q��������U����?  |f�E�f��f�E��M�Q�U�R�ƾ�����Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�K�������}� },�E���%�   �E��	�M����M��}� ~�U�R�.�������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P�֫�����M�Q�ʫ�����U�R�E�P�ʠ�����M�Q讫�����U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�R�E�Q�`������E��}� t0�U��Rj�E�HQ�?������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�
������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR�ի������]�������������������������������������������������̋�U��j
j �EP�ˢ����]���������̋�U��EPj
j �MQ襤����]���������������������̋�U��EP������]�������������̋�U��EP�MQ������]���������̋�U��j
j �EP臜����]���������̋�U��EPj
j �MQ�O�����]����������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� �������������������������������������������U��SVWUj j h��
�u臫��]_^[��]ËL$�A   �   t2�D$�H�3��d���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��
d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��
u�Q�R9Qu�   �SQ�P��SQ�P��L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������������������̋�U���8�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh�j jphj�b�������u̃}� u.�����    j jphhX{h�����������   3Ƀ} ���MЃ}� uh�<j juhj���������u̃}� u.豹���    j juhhX{h�<贱��������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P�������E��} u�E��Q�M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �p������EȋE���]������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�l�����]�������������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h�j h�  hj�/�������u̃}� u.�����    j h�  hht{h�����������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQhA9������]������������������̋�U��EP�MQ�URhA9�١����]����������������̋�U��EPj �MQh=諡����]������������������̋�U��EP�MQ�URh=�y�����]����������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh�j jphj�b�������u̃}� u.�����    j jphh�{h�����������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh�j jshj��������u̃}� u.蛵���    j jshh�{h�螭���������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �C������Eă}��t�E���UU�B� �E��x }�����������]��������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPhA9�������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhA9蹸�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�|j h�   hj�\�������u̃}� u1�����    j h�   hh\|h�|�����������  �} t�} v	�E�   ��E�    �U�U�}� u!h|j h�   hj�ܒ������u̃}� u1菲���    j h�   hh\|h|菪��������d  �MQ�UR�EP�MQ�URh<�h������E��}� }U�E�  �}�tI�}���t@�}v:�M��9<�s�<��U��	�E���E�M�Qh�   �U��R��������}��uu3�t	�E�   ��E�    �M�M��}� u!h�{j h�   hj�ߑ������u̃}� u.蒱��� "   j h�   hh\|h�{蒩��������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9<�s
�<��E���M����U+щU��E�Ph�   �M��U�D
P�������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�5�����]���������������̋�U���,�E������E�    3��} ���E�}� u!h�|j h  hj�%�������u̃}� u1�د���    j h  hh�|h�|�ا��������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!h|j h  hj茏������u̃}� u1�?����    j h  hh�|h|�?���������|  �M;M��   ������U��EP�MQ�UR�E��P�MQh<��������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9<�s�<��U���E���M+ȉM�U�Rh�   �E�M�TR膏�����i����8"u
�_����M������  �`�K�����U��EP�MQ�UR�EP�MQh<�K������E��UU�B� �}��u"�}�u�����8"u
������M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U��E�Ph�   �M��Q詎�����}��uu3�t	�E�   ��E�    �E܉E�}� u!h�{j hB  hj茍������u̃}� u.�?���� "   j hB  hh�|h�{�?�������������z�}�t\�}���tS�U���;UsH�E����M+�9<�s�<��U���E����M+ȉM؋U�Rh�   �E��M�TR�Ǎ�����}� }	�E�������E��EԋEԋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�Y�����]�����������̋�U����EPj �MQ�UR�EPh=�{������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh=�������E��}� }	�E�������U��U��E���]������������������������̋�U��j�hH�h)d�    P���SVW���1E�3�P�E�d�    �E������E������}�u!藓���     �f���� 	   ��������  �} |�E;�s	�E�   ��E�    �MԉM܃}� uh@~j jMh�}j�L�������u̃}� u<�%����     ������ 	   j jMh�}h�}h@~��������������C  �E���M������@�D
������؉E�uh|}j jNh�}j�É������u̃}� u<蜒���     �k���� 	   j jNh�}h�}h|}�n������������   �UR�������E�    �E���M������@�D
��t �MQ�UR�EP�MQ�a������E��U��F����� 	   �����     �E������E�����3�uh�|j jYh�}j��������u��E������   ��MQ�m�����ËE��U�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��UR�ѕ�����E�}��u;讧��� 	   3�u!h�|j h�   h�}j�Ň������u̃������   �UR�E�P�M�Q�U�R��"�E��}��u#�$"�E��}� t�E�P�������������>�M���U������@�L����U���E������@�L�E��U���]������������������������������������������������������������������������̋�U��j�hh�h)d�    P���SVW���1E�3�P�E�d�    �}�u蕏���     �d���� 	   ����  �} |�E;�s	�E�   ��E�    �M؉M��}� uh@~j jCh�~j�M�������u̃}� u9�&����     ������ 	   j jCh�~h�~h@~�����������/  �E���M������@�D
������؉E�uh|}j jDh�~j�ǅ������u̃}� u9蠎���     �o���� 	   j jDh�~h�~h|}�r���������   �UR�������E�    �E���M������@�D
��t�MQ�UR�EP踀�����E��?������ 	   �����     �E�����3�uh�|j jOh�~j���������u��E������   ��EP肀����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U�츐<  蹂�����3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uh�j jmh�~j�̓������u̃}� u9覌���     �u����    j jmh�~h�h��x���������
  �E���M������@�D
$�����E��M���t	�U���uo�E��������E�uhtj juh�~j�+�������u̃}� u9�����     �Ӣ���    j juh�~h�ht�֚���������	  �U���E������@�T�� tjj j �EP�������MQ芛������td�U���E������@�T��   tA������EԋEԋHl3҃y �U�E�P�M���U������@�Q��"�E�}� ��  �}� t�U�����  ��"�E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M������@�|
8 ��   �E���M������@�D
4P�{������u!h0j h�   h�~j�w�������u̋U���E������@�T4�U��EЊ�M��U���E������@�D8    j�U�R�E�P�Y��������u�  �   �M��R�"{��������   �E�+E�M+ȃ�v'j�U�R�E�P���������u�O  �MЃ��M��K�U���E������@�UЊ�T4�E���M������@�D
8   �E����E���  �j�M�Q�U�R��������u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R��!�Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M������@�
P��"��t�M�+MM�M��U�;U�}�  ��$"�E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M������@�
P��"��t!�M�;M�}�   �U���U�E����E���$"�E��   �   �M���t	�U���u{�E�P�[��������U�;�u�E����E���$"�E��R�}� tG�E�   �   f�M��U�R���������M�;�u�U����U��E���E���$"�E���t�����  �M���U������@�L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E������@�R��"��t �E�E��E�������������+�9M�}���$"�E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U������@�Q��"��t �U�U��U�������������+�9E�}���$"�E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  ��!��t�����t��� u�$"�E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E������@�R��"��t��p���E���p�����$"�E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U������@�Q��"��t�E�    �U��U��	�$"�E�}� ��   �}� t0�}�u�C���� 	   �^����M���U�R��v��������V�L�E���M������@�D
��@t�M���u3��%������    �����     ������E�+E�M�3��X�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} uh�Aj j.h �j�v������u̋X����X��U�U�j:h�jh   �o�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������������������������������������������������������̋�U����}�u�ٔ��� 	   3��   �} |�E;�s	�E�   ��E�    �M��M��}� uh@~j j(h��j��t������u̃}� u*�v���� 	   j j(h��h��h@~�y�����3���E���M������@�D
��@��]���������������������������������������������������̋�U��h�]����̋�U��Q�=� u��   ��=�}
��   h�   h$�jj��P諒�����l��=l� u?��   h�   h$�jj��Q�v������l��=l� u
�   �   �E�    �	�U����U��}�}�E���h��M��l������E�    �	�E����E��}�}f�M����U�������@�<�t8�M����U�������@�<�t�M����U�������@�< u�M���ǁx������3���]������������������������������������������������������������������������������������̋�U���,v�������t��x��j�l�Q轅����]�������������������̋�U��}h�r4�}��w+�E-h�����P��s�����M�Q�� �  �E�P��M�� Q��"]�������������������������������̋�U��}}#�E��P�ls�����M�Q�� �  �E�P��M�� Q��"]�������������������̋�U��}h�r4�}��w+�E�H������U�J�E-h�����P��������M�� Q��"]�������������������������������̋�U��}}#�E�H������U�J�E��P艃������M�� Q��"]�������������������̋�U��Q3��} ���E��}� uh�Dj j)hp�j�p������u̃}� u+�K����    j j)hp�h\�h�D�N����������U�B��]�������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    3��} ���E؃}� uh�j j6h��j��o������u̃}� u.菏���    j j6h��h�h�蒇��������   �U�U��Ā���� Pj�ڑ�����E�    誀���� P��n�����E܋E�Pj �MQ茀���� P迀�����E��x����� P�U�R�Ӌ�����E������   ��U����� Pj������ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP��g������]������������̋�U��Q�E�E��M�Q�UR�EP�u������]������������̋�U��Q�E�E��M�Qj �UR�u������]��������������̋�U��Q�E�E��M�Q�UR�EP�_u������]������������̋�U��Q�E�E��M�Qj �UR�1u������]��������������̋�U��������3�9\����M��} t������U���E�    �E��\��E���]������������������������̋�U������3�9\�����]��������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh��j jJh��j��l������u̃}� u0�x����    j jJh��hl�h���{������   �\  �UR�M��:z���M���k��� �x ��   �M���   ~C�} t�} v�URj �EP�m���������� *   ������M؍M�轌���E���  �} tw3�;U��؉E�uhd�j j]h��j��k������u̃}� u=衋��� "   j j]h��hl�hd�褃�����E�"   �M��H����E��x  �U�E��} t	�M�   �E�    �M������E��J  �=  �E�    �U�Rj �EP�MQj�URj �M��j��� �HQ��!�E��}� t
�}� ��   �}� ��   �$"��z��   �} t�} v�URj �EP��k����3�t	�E�   ��E�    �U��U܃}� uh�{j j{h��j�j������u̃}� u:�r���� "   j j{h��hl�h�{�u������E�"   �M������E��L�8���� *   �-�����MȍM�������E��*�} t�U�E���E�    �M��Պ���E���M��Ȋ����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�zs����]��������������̋�U��� �E������EP�M���v���M��ch��P�MQ�M��Uh������   P�MQ�U�R� s�����E�}� u�E��E���E������M��M�M��c����E��]�����������������������������������������̋�U����E�����j �EP����P�MQ�U�R�r�����E��}� u�E��E���E������E��]���������������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uh��j jEhh�j��g������u̃}� u.苇���    j jEhh�h4�h�����������  �MQ�M��Ou���} �  �M���f����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M�������E��O  �M����M��U���U뱋E��EԍM�趇���E��%  �  �MQ�URj��EPj	�M��Df����QR��!�E��}� t�E����EЍM��k����E���  �$"��zt*�|���� *   3ɋUf�
�E������M��6����E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M��e��P�M��R�/h������t@�E��H��u,������ *   3ҋEf��E������M�贆���E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M��,e����QR��!�E��}� u*舅��� *   3��Mf��E������M��B����E��   �U��U��M��,����E��   �   �M���d��� �x u�MQ�i�����E��M�������E��j�`j j j��URj	�M��d��� �HQ��!�E��}� u!����� *   �E������M�讅���E�� ��U����U��M�薅���E���M�艅����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�UR�EP�ol����]�����������������̋�U��=L� uh��EP�MQ�UR�ʆ������j �EP�MQ�UR谆����]�����������������������������̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!h��j h�   hh�j�c������u̃}� u3�͂���    j h�   hh�hd�h����z�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���E��M���Qh�   �U��R�Xc�����} t	�E�     �MQ�M��p���U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h0�j h  hh�j�b������u̃}� u@�ˁ���    j h  hh�hd�h0���y�����E�   �M��o����E���  �M��a��P�E�P�MQ�UR�3j�����E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���M��U���Rh�   �E��P�$b����������MЍM��с���E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9<�s�<��M��	�U���U��E���Ph�   �M��Q�a�����U�9U����E�u!h��j h  hh�j�`������u̃}� u=�4���� "   j h  hh�hd�h���4x�����E�"   �M��؀���E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM�蝀���Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�p����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�.j jhXGj�^������u̃}� u0�S~���    j jhXGh4�h�.�Vv�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U��E�Ph�   �M��Q��^����3҃} �U��}� uh�-j jhXGj��]������u̃}� u0�}���    j jhXGh4�h�-�u�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9<�s
�<��E��	�M���M܋U�Rh�   �E��P��]������F��t3�t	�E�   ��E�    �E؉E�}� uh�Fj j hXGj��\������u̃}� u0�|���    j j hXGh4�h�F�t�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9<�s
�<��E��	�M���MԋU�Rh�   �E��P��\������-��t3�t	�E�   ��E�    �EЉE�}� uh<-j j*hXGj��[������u̃}� u-�u{��� "   j j*hXGh4�h<-�xs�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9<�s�<��U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR��[����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uh,�j jfhX�j�vY������u̃}� u0�)y���    j jfhX�hH�h,��,q�����   ��  3�;U��؉E�uh �j jghX�j�Y������u̃}� u0��x���    j jghX�hH�h ���p�����   �  �U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���UԋE�Ph�   �M��Q�_Y����3҃} ��;U��؉E�uh��j jihX�j�SX������u̃}� u0�x��� "   j jihX�hH�h���	p�����"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uh��j jjhX�j��W������u̃}� u0�w���    j jjhX�hH�h���o�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!hL�j h�   hX�j��V������u̃}� u0�v��� "   j h�   hX�hH�hL��n�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ������]�����������������̋�U��j �EP�MQ�UR�EP�T���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!h,�j h>  hX�j�MT������u̃}� u3� t���    j h>  hX�hȆh,�� l�����   �,  3�;U���؉E�u!h �j h?  hX�j��S������u̃}� u3�s���    j h?  hX�hȆh ��k�����   ��  �U�� �}��tI�}����t@�}�v:�EЃ�9<�s�<��M��	�UЃ��ŰE�Ph�   �Mԃ�Q�-T����3҃} ��;U���؉E�u!h��j hA  hX�j�S������u̃}� u3��r��� "   j hA  hX�hȆh����j�����"   ��  �}r�}$w	�E�   ��E�    �UȉU܃}� u!h��j hB  hX�j�R������u̃}� u3�Or���    j hB  hX�hȆh���Oj�����   �{  �E�    �MԉM��} t+�U��-�E����E��M����M��U�ڋE�� �؉U�E�M��M�U3�PR�MQ�UR�r���E�E3�QP�UR�EP�1p���E�U�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} w�} v�U�;U�r��E�;E�rl�M�� �U�;U���؉E�u!hL�j hf  hX�j�cQ������u̃}� u0�q��� "   j hf  hX�hȆhL��i�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�B���]����������������̋�U���x���3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uh��j jfh�j�[O������u̃}� u.�o���    j jfh�h��h���g��������8  �UR�M���\���} �.  �M��QN��� �x ��   �M�;Msp�U�=�   ~"�n��� *   �E������M��co���E���  �MM��U���M��E���E��u�M��M��M��-o���E��  �U����U�눋E��E��M��o���E��  �  �M��M������   ��   �} v�UR�EP�  ���E�M�Qj �UR�EP�MQ�URj �M��bM��� �HQ��!�E��}� t3�}� u-�UU��B���u	�M����M��U��U��M��on���E���  �m��� *   �E������M��Mn���E���  ��  �E�Pj �MQ�URj��EPj �M���L����QR��!�E��}� t�}� u�E����E��M���m���E��j  �}� u�$"��zt"�m��� *   �E������M���m���E��7  �M�;M�  �U�Rj �M��TL��� ���   Q�U�Rj�EPj �M��7L����QR��!�E�}� t�}� t"�l��� *   �E������M��Om���E���  �}� |�}�v"�_l��� *   �E������M��!m���E��  �E�E�;Ev�M��M��M�� m���E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M��l���E��  벋U���U������E��E��M��l���E���   ��   �M��#K����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"�\k��� *   �E������M��l���E��   �Ũ��U�벋ẺE��M���k���E��t�j�M�Qj j j j��URj �M��J��� �HQ��!�E��}� t�}� t��j��� *   �E������M��k���E���U����U��M��k���E���M��k���M�3��;n����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�������������������������������������̋�U��EP�MQ�UR�EP�c����]�����������������̋�U��j �EP�MQ�UR�vc����]�������������������̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h �j h@  h�j�ZH������u̃}� u3�h���    j h@  h�h܇h ��`�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U��E�Ph�   �M��Q�H�����} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h0�j hL  h�j�hG������u̃}� u3�g���    j hL  h�h܇h0��_�����   �  �MQ�U�R�EP�MQ�a�����E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9<�s�<��M��	�U���U؋E�Ph�   �M��Q�G�����lf��� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9<�s
�<��E��	�M���MԋU�Rh�   �E��P� G�����M9M���ډU�u!h��j hd  h�j��E������u̃}� u0�e��� "   j hd  h�h܇h���]�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ��D����]�����������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h�j h�   h؈j�?D������u̃}� u1��c���    j h�   h؈h��h���[��������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h�j h�   h؈j�C������u̃}� u1�rc���    j h�   h؈h��h��r[��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �[�����Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj �Z�����E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh�H�O�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh�H� O�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�|j h  h؈j�@������u̃}� u1�_`���    j h  h؈h��h�|�_X���������  �} t�} v	�E�   ��E�    �U�U�}� u!hP�j h  h؈j�,@������u̃}� u1��_���    j h  h؈h��hP���W��������j  �MQ�UR�EP�MQ�URh�8��M�����E��}� }X3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���M�U���Rh�   �E��P�I@�����}��uu3�t	�E�   ��E�    �U�U��}� u!h�{j h  h؈j�,?������u̃}� u.��^��� "   j h  h؈h��h�{��V��������m�}� |d�}�t^�}���tU�M���;MsJ�U����E+�9<�s�<��M���U����E+E��M���Qh�   �U��E�LPQ�d?�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�H����]���������������̋�U���,�E������E�    3��} ���E�}� u!h�|j h9  h؈j�u=������u̃}� u1�(]���    j h9  h؈hȉh�|�(U��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!hP�j h?  h؈j��<������u̃}� u1�\���    j h?  h؈hȉhP��T��������  �M;M��   �R\����U��EP�MQ�UR�E��P�MQh�8�fJ�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9<�s�<��U���E���M+ȉM�U���Rh�   �E�M�TAR��<�����[���8"u
�[���M�������  �c�[����U��EP�MQ�UR�EP�MQh�8�I�����E�3ҋE�Mf�TA��}��u"�}�u�N[���8"u
�D[���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9<�s
�<��E��	�M���M��U���Rh�   �E��P��;�����}��ux3�t	�E�   ��E�    �U܉U�}� u!h�{j hf  h؈j��:������u̃}� u1�Z��� "   j hf  h؈hȉh�{�R��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9<�s�<��M���U����E+E؋M���Qh�   �U��E�LPQ�;�����}� }	�E�������U��UԋEԋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�H����]�����������̋�U����EPj �MQ�UR�EPhn9��F�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhn9�`F�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uh,�j jfhX�j�7������u̃}� u0�9W���    j jfhX�h��h,��<O�����   �  3�;U��؉E�uh �j jghX�j�$7������u̃}� u0��V���    j jghX�h��h ���N�����   �  3ҋEf��}�tK�}���tB�}v<�M��9<�s�<��U��	�E���EԋM���Qh�   �U��R�k7����3��} ����;E��ىM�uh��j jihX�j�_6������u̃}� u0�V��� "   j jihX�h��h���N�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uh��j jjhX�j��5������u̃}� u0�U���    j jjhX�h��h���M�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!hL�j h�   hX�j��4������u̃}� u0�T��� "   j h�   hX�h��hL��L�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�e�����]�����������������̋�U��j �EP�MQ�UR�EP�4���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!h,�j h>  hX�j�=2������u̃}� u3��Q���    j h>  hX�h �h,���I�����   �A  3�;U���؉E�u!h �j h?  hX�j��1������u̃}� u3�Q���    j h?  hX�h �h ��I�����   ��  3ҋE�f��}��tK�}����tB�}�v<�MЃ�9<�s�<��U��	�EЃ��E̋M���Qh�   �Uԃ�R�2����3��} ����;E���ىM�u!h��j hA  hX�j�
1������u̃}� u3�P��� "   j hA  hX�h �h���H�����"   �  �}r�}$w	�E�   ��E�    �EȉE܃}� u!h��j hB  hX�j�0������u̃}� u3�;P���    j hB  hX�h �h���;H�����   �  �E�    �UԉU��} t0�-   �M�f��U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ��O���E�U3�PR�MQ�UR�N���E�U�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} w�} v�M�;M�r��U�;U�rn3��M�f��U�;U���؉E�u!hL�j hf  hX�j�F/������u̃}� u0��N��� "   j hf  hX�h �hL���F�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�"���]����������������̋�U����  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���:���E�    ��L���E�3Ƀ} �������������� u!h�Dj h  h�Dj��,������u̃����� uF�L���    j h  h�Dh�h�D�D����ǅ<��������M��BM����<����  3��} �������������� u!h�j h  h�Dj�i,������u̃����� uF�L���    j h  h�Dh�h��D����ǅ8��������M��L����8����!  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U����  ������ ��  �������� |%��������x���������A����,����
ǅ,���    ��,������������������������B����������������(�����(����*  ��(����$��	�E�   ������Q�UR������P�h  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ��������$�����$����� ��$�����$���wL��$�����,
�$�
�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�4G�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP��F�����Ẽ}� }�E�������M�k�
�������DЉE��  �������� ����� �����I�� ����� ���.�  �� �����T
�$�@
�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  ��������
�$��
�M���0  u	�U��� �U��E�   �EP�E����f�������M��� tW���������   ������ƅ���� �M��A'��P�M��8'��� ���   Q������R������P�E������}�E�   �f������f�������������U��E�   �  �EP�|D���������������� t�������y u�`��U��E�P�+�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ����������������MQ�C�����E��U��� ��   �}� u�`��E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M��%��P�������Q�9(������t������������������������������d�}� u	�d��M��E�   �U���|�������������������������t��|������t��|�������|����ɋ�|���+U����U��  �EP�B������x����6������   3�tǅ���   �
ǅ���    �������t�����t��� u!h�Bj h�  h�Dj�\%������u̃�t��� uF�E���    j h�  h�Dh�h�B�=����ǅ4��������M��E����4����  ��  �M��� t��x���f������f����x�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  htBj�Ḿ�]  Q������E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��A#��P�U�R�E�P������Q�U�R�E�P��h���Q��R��!�Ѓ��E�%�   t%�}� u�M���"��P�M�Q��R��!�Ѓ���������gu)�M���   u�M���"��P�U�R��P��!�Ѓ��M����-u�E�   �E��M����M��U�R�o'�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�+������X�����\����   �U���   t�EP�p+������X�����\����   �M��� tB�U���@t�EP�%?��������X�����\�����MQ�	?���������X�����\����=�U���@t�EP��>�������X�����\�����MQ��>����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R��@����0��d����E��RP��T���P��P���Q��>����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �]  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��>��P�M��5������   R��H���P������Q�<������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��L���Rj �  ���}� tj�E�P�y1�����E�    �"�����������0����M��>����0����M�3��EA����]Ð��
��
�
y�
��
��
�
P�
R�
]�
G�
<�
k�
t�
 �I ��
4�
R�
?�
K�
 �
��
� �= "��
��� ���   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ��0�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U���@�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h�j h�   h؈j�������u̃}� u1�R6���    j h�   h؈h4�h��R.��������V  3Ƀ} ���MЃ}� u!h�<j h�   h؈j�5������u̃}� u1��5���    j h�   h؈h4�h�<��-���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P�6�����E��} u�E��   �M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �-�����EȋE��H���MċU��EĉB�}� |!�M��� 3�%�   �E��M�����E����M�Qj �T-�����E��E���]��������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�0����]�������������������̋�U��EP�MQ�UR�EP��/����]�����������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h�j h�  h؈j��������u̃}� u.�3���    j h�  h؈hT�h��+��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh�H�)����]������������������̋�U��EP�MQ�URh�H�T)����]����������������̋�U��EPj �MQhn9�&)����]������������������̋�U��EP�MQ�URhn9��(����]����������������̋�U���@���3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �M�y ��  �U�z u+�E��Ph  �M�Q0Rj �E�P�3������t�"  j^h@�jj������E�jbh@�jjh�  �t0�����E�jdh@�jjh�  �Y0�����E�jfh@�jjh�  �>0�����E�jhh@�jjh  �#0�����E�}� t�}� t�}� t�}� t�}� u�}  �M��    �U�U��E�    �	�E����E��}�   }�M��U���E����E��ۍM�Q�U�BP��"��u�&  �}�v�  �M܉Mă}�~S�U�U��	�E����E��M����t8�E��H��t-�U���E��	�M����M��U��B9E��M�M�� ���j j �U�BP�Ḿ�   Qh   �U�Rjj �8!���� ��u�  j �E�HQh�   �Uȁ   Rh�   �E��Ph   �M�QRj �0"����$��u�E  j �E�HQh�   �U��   Rh�   �E��Ph   �M�QRj ��!����$��u�  3��M�f���   �U��B �E��@ �M�Ɓ�    �U�Ƃ�    �}�~]�E�E��	�M����M��U����tB�M��Q��t7�E���M��	�U����U��E��H9M�� �  �E��M�f��A   ���h�   �Ú�   R�E�P�$����j�Mȁ�   Q�U�R�����j�E�   P�M�Q�������U���    ��   �E���   Q�("����   3�uj j h�   hȊj�������u�j�M���   ���   R��!����j�E���   ��   Q�!����j�U���   -�   P�!����j�M���   R�!�����E��    �M�UЉ��   �E�   �M���   �Ú��   �E���   �Mȁ��   �U���   �E��   �M���   �U�Eĉ��   j�M�Q�!����3���   j�U�R�!����j�E�P�� ����j�M�Q�� ����j�U�R�� ����j�E�P�� �����   �   �   �M���    tA�U���   P�("��u-�M���    w!h��j h�   hȊj�������u̋Eǀ�       �Mǁ�       ��o�E���   �(t�U���   ��u�M���   �Uǂ�      3��M�3��0����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�������E��E��Hl�M��U�;�t�E��Hp#H�u�g���E��U����   ��]�������������������������̋�U��Q�} u
�R'���E���E����   �U��E���]���������������������̋�U�������E��E��Hl�M��U�;�t�E��Hp#H�u�����E��U��B��]����������������������������̋�U�������E��E��Hl�M��U�;�t�E��Hp#H�u�g���E��U��B��]����������������������������̋�U����D���E��E��Hl�M��U�;�t�E��Hp#H�u����E��E�����]����������������������������̋�U��3�]��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^���������������������������̋�U��Q�E�    �} u3��S  �}��   �	�E����E��M��9M���   �U���U�E���E�M�Q���t�E�H��U�B�;�t�M�A��U�J�+���   �U�B���t�M�Q��E�H�;�t�U�B��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��X�����	�E����E��M�;Ms>�U���t�M��E�;�t�U��M�+���E���E�M���M�3���]������������������������������������������������������������������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U���(�E�E��M�M��U�U��}��g  �E��$��"�M�Q�U�R��  ���E�}� t�E�E��s�M���Q�U���R��  ���E�}� t�E�E��F�M���Q�U���R�  ���E�}� t�E�E���M���Q�U���R�  ���E�E�E�M�M�E���   �U�R�E�P�Y  ���E�}� t�M�M��F�U���R�E���P�2  ���E�}� t�M�M���U���R�E���P�  ���E܋M܉M��E��i�U�R�E�P��   ���E�}� t�M�M���U���R�E���P��   ���E؋E��*�M�Q�U�R�   ���3���EP�M�Q�U�R�  ����]Ðw"e"&"�!!�����������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��+�P�   ����]�����������������̋�U��} t3��} ���D ��E�E]����������������̋�U����} �R  �EP�MQ�Q	  ���E��}� t�E��O  �U��R�E��P�*	  ���E��}� t�E��(  �M��Q�U��R�	  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�g  ���E��}� t�E��e  �U��R�E��P�@  ���E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$�*�U��R�E��P��  ���E��}� t�E���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��}  �U��R�E��P�X  ���E��}� t�E��V  �M��Q�U��R�1  ���E��}� t�E��/  �E��P�M��Q�
  ���E��}� t�E��  �U��R�E��P��  ���E��}� t�E���  3���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��  �U��R�E��P�g  ���E��}� t�E��e  �M��Q�U��R�@  ���E��}� t�E��>  �E��P�M��Q�  ���E��}� t�E��  �U��	R�E��	P��  ���E��}� t�E���  �M��Q�U��R��  ���E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�b  ���E��}� t�E��`  �E��P�M��Q�;  ���E��}� t�E��9  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���E��}� t�E���  �E��
P�M��
Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���  �E��P�M��Q�]  ���E��}� t�E��[  �U��R�E��P�6  ���E��}� t�E��4  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���   �U��R�E��P��  ���E��}� t�E��   �M��Q�U��R�  ���E��}� t�E��   �E��P�M��Q�s  ���E��}� t�E��t�U��R�E��P�o������E��}� t�M��M��F�U��R�E��P�H������E��}� t�M��M���U��R�E��P�!������E��M��M�E��3���]Ë�1&I'u(�)
&"'N(z)�%�&'(S)�%�& (,)�%�&�')n%�&�'�(G%_&�'�( %8&d'�(�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��;�tK�E�E��M�M�U�R�E�P�������E�}� t�M�M���U���R�E��P�\������E�E��3���]�������������������������������������������̋�U��� �E�E��M�M��U��E��
;��   �U�U��E�E�M�Q�U�R��������E�}� t�E�E��s�M���Q�U��R�������E�}� t�E�E��F�M���Q�U��R�������E�}� t�E�E���M���Q�U��R�n������E��E��E�M�M�E��3���]�����������������������������������������������������������������̋�U����4���   �E��} u�E�P�\  ���  �M��U��E��@�M��A�U��z t#�E��H���t�E���Pjh����  ���M��A    �U��: ��   �E�������   �E��x t�M��Q���t�M�Q�O  ����U�R�	  ���E��x uG�M�Qj@hP��u  ����t0�U��z t�E��H���t�E�P��  ����M�Q�1	  ���0�U��z t�E��H���t�E�P�  ����M�Q�?  ���U��z u3��N  �} t�E�   �E���E�    �M�Q�U�R�U  ���E��}� t!�}���  t�}���  t�E�P��"��u3���   j�M��QR� #��u3���   �} t&�E�M�f�Qf��E�M�f�Qf�P�Ef�M�f�H�} ��   �U�=  u4j h1  h(�h�hДh��j@�MQ�����P�]����� j@�URh  �E��HQ��"��u3��Bj@�U��@Rh  �E��HQ��"��u3��j
j�U�   R�E�P�������   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�;Eb�}� t\�E�E�+����E��M��U��P�M�R������E�}� u�E��M�T��E���}� }�M����M�	�U����U��3��}� ����]�����������������������������������̋�U��Q�E�Q�������3҃��E�P�M�QR�������3Ƀ����U�J�E�@    �M�y t	�E�   ��U�P��  ���E��M�U��Qjh 3�#�E�H��   t�U�B%   t�M�Q��u
�E�@    ��]����������������������������������������������������������̋�U���   ���3ŉE��7 ���   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q��"��u��|����B    �   �  �E�P��|����QR���������r  jx�E�P��|����Q��ҁ������  R��x���P��"��u��|����A    �   �G  �U�R��|����Q�\������u:��|����B  ��|����A��|�����x����B��|�����x����Q��   ��|����H����   ��|����z tt��|����HQ�U�R��|����Q�B������uQ��|����B����|����A��|�����x����B��|����R�i�������|���;Au��|�����x����B�E��|����Q��u7��x���P��  ����t$��|����Q����|����P��|�����x����Q��|����H��   ��   ��  jx�U�R��|����H��Ɂ������  Q��x���R��"��u��|����@    �   �  �M�Q��|����P���������
  ��|����Q��   ��|����P��|����y t7��|����B   ��|����A��|����z u��|�����x����H�   ��|����z tl��|����Q��������|���;BuP��|���Pj��x���Q��  ����t2��|����B   ��|����A��|����z u��|�����x����H�2��|����B   ��|����A��|����z u��|�����x����H�   ��|����z ut��|����x th�M�Q��|����P�������uO��|���Qj ��x���R�C  ����t3��|����H��   ��|����J��|����x u��|�����x����Q��|����@��������M�3�� ����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�Q������3҃��E�P�M�y t	�E�   ��U�P��  ���E��M�U��Qjh�8�#�E�H��u
�U�B    ��]��������������������������������������������̋�U���   ���3ŉE��G����   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q��"��u��|����B    �   �  �E�P��|����R��������u`��|����x u��|���Qj��x���R�y  ����t3��|�����x����H��|�����x����B��|����Q����|����P�   ��|����y ut��|����z th�E�P��|����R�A������uO��|���Pj ��x���Q��  ����t3��|�����x����B��|�����x����Q��|����H����|����J��|����@��������M�3������]� ������������������������������������������������������������������������������������������������������̋�U��E�HQ������3҃��E�PjhP;�#�M�Q��u
�E�@    ]��������������������������̋�U���   ���3ŉE�������   ��|����EP�B  ����x���jx�M�Q��|����B���%���  P��x���Q��"��u��|����B    �   �s�E�P��|����QR�t������uF��x���P��  ����t3��|�����x����Q��|�����x����H��|����B����|����A��|����B��������M�3�������]� ������������������������������������������������������������������̋�U��Q�E�H��  �U�J�#�E��E�M��H�U�E��B��]�������������������������̋�U��Q�} t�E���th���UR�T�������u0j�E�Ph  �M�QR��"��u3��Y�}� u��"�K�Fh���EP��������u"j�M�Qh   �U�BP��"��u3����MQ�|	�����E��E���]��������������������������������������������������������̋�U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E��;�u3���ظ   ��]����������������������̋�U���V�E%�  �ȁ�   �щU�j�E�Ph   �M�Q��"��u3��9�U;U�t,�} t&�E�Q��   �����U�P������;�u3���   ^��]������������������������������������̋�U����E�    �E��M��U��E���E��tM�M���a|�U���f�E���'�E���M���A|�U���F
�E����E��M����U��DЉE�뚋E���]������������������������������������̋�U����E�    �E��M��U���U�E���A|	�M���Z~�U���a|%�E���z�M����M��U��E��M���M���E���]�������������������������̋�U���EP�MQ�s�����]�������̋�U��Q�E=��  u3��G�M��   }�U���P�M#��&�U�Rj�EPj��"��u3�f�M��E��U#�]��������������������������������̋�U���EP�MQ�������]�������̋�U���������   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR�������   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�i   �� �   ��]���������������������������������������������������������������������������������������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}��
����E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  �T������    u��  �A������   �E�3������   �M�E�j�UR���������t��m����E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u�'�����������    ty�������   �E�����ǀ�       �M�Q�UR��  ������t�C�M�Q�  ���Ѕ�t+j�EP�7�����h���M������h���M�Q�����������U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP��������E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q��������u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�  ��,�	���D���������M��tj�UR�������E�����   �M��������!���   �E�x ��   �M�QR�EP��  ���ȅ���   �[������   �U��M������   �E��?����M���   �1����U���   �}$ u�EP�MQ�������UR�E$P�����j��MQ�UR�EP�_������M�QR�C  ��������M���   ������U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP�  �� ��T����~������    u��������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M��EP�M��B����M�����E���]� ��������̋�U��Q�M��E�� ���M��A ����]������������������̋�U��Q�M��M��b����E��t�M�Q�s������E���]� �����������������̋�U��Q�M��EP�M�������M�����E���]� ��������̋�U���V�E�8  �u�c  �S������    tW�E����������9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP��������t��   �M�y t��C����U�R�E�P�MQ�U R�EP��������E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������������������������������������������������������������������������������������������������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�:�������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����������������������������������������������������̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@�g���ǀ�       �)����S������    ~�E����   �E�M����E�3��3���]�������������������������������������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E������   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}������M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R�����E�    ��E�P������Ëe��E�    �M��M��f����E������   �)��������    ~������   �EԋUԋ���MԉËU�;Uu�������E�M�H�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����E�E��}  t�M Q�UR�E�P�MQ��������}, u�UR�EP������MQ�U,R�����E$�Q�UR�EP�M�Q�(������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�T   ���E��}� t�EP�M�Q������]�������������������������������������������������������̋�U��j�h@�h)d�    P���SVW���1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R�������E���������   �E��������   �M������U���   �����M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP�G������E��E�    ��   �M�Q�N  ��Ëe��C���ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP��������E�    �E�    �E������E�    �   �   �M�U��Q��E�P�t������?����Mȉ��   �1����Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP��������t�M�Q�UR������ËEЋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u����ǀ     �   ��3���]�����������������������������������̋�U��j�hp�h)d�    P���SVW���1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR��������t9j�E�P�{�������t'�M��U�B��M��Q�U��P�~������M���������@  �U���txj�M�QR�9�������tYj�E�P��������tG�M�QR�E�HQ�U�R�������E�xu"�M��9 t�U��R�E��Q��������U����W����   �E�x uZj�M�QR��������t>j�E�P��������t,�M�QR�E��P�M�QR������P�E�P�r������������[j�M�QR�^�������tAj�E�P�>�������t/�M�QR��������t�E���t	�E�   ��E�   ������E�������   Ëe�������E������E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�.������E��}�t�}�t+�R�U��R�E�HQ������P�U�BP�M�Q�P����)j�U��R�E�HQ������P�U�BP�M�Q������E�������   Ëe��?����E������M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h��h)d�    P��SVW���1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR������E�������E�����Ëe��L����E������M�d�    Y_^[��]�������������������������������������������������̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]������������������������̋�U�������3Ƀ��    ����]������̋�U���(�} u3���  �E��M��} t�U�B����   �M��9MOC�t�U��:RCC�t�E��@uz�M��9csm�uK�U��zuB�E��x �t�M��y!�t�U��z"�u�E��x u�������    u3��I  �����   �E܋M܋���E܉�   �%  �M��9csm��  �U��z�  �E��x �t�M��y!�t�U��z"���   �E��x u#�������    u3���   �������   �M��U�U�E�E��M���   ��M��U��B�H���M�U��B�H��U���E����E��M���M�}� ~d�U��E��M��QR�E�P�M�Q���������t?� ����   �E؋U؋���M؉�} t�U�R�E�P�MQ�U�R�������   ��3���]�����������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E��M����M�U���U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u�������   �E��M��QR�E�P�^������E������M􋐈   ������M����   ��r����M����   ��U�������E�� �����P����   �E�M����E��6������    }�(���ǀ�       �   ��]������������������������������������������������������������������������������������̋�U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!�a����   �E��U�����M���   �3���]����������������������������������������������̋�U����E�E��M����M�U���U��E�8��G  �M�Q�	������} ��   ��������   �:csm�u~�������   �xum�������   �y �t(�������   �z!�t�~������   �x"�u1�j������   �QR��������tj�M������   P�������9������   �9csm�um�&������   �zu\�������   �x �t(�������   �y!�t��������   �z"�u �} t������   �E��E�����U��
�����M����   �����M�����   ��]���������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U��j�h��h)d�    P��SVW���1E�3�P�E�d�    �e��E�    �M�U�E�������E�P�\�����Ëe��E������M�d�    Y_^[��]��������������������������������������������̋�U��j�h��h)d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�U���E�������M�Q������Ëe��E������M�d�    Y_^[��]����������������������������������������̋�U��j�h�h)d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�U�E�������M�Q������Ëe��E������M�d�    Y_^[��]�������������������������������������������̋�U��j�h0�h)d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�MQ�UR�EP�U�E�������M�Q�o�����Ëe��E������M�d�    Y_^[��]�����������������������������������������������̋�U����} t�������} u�B����E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR���������t�E���뀊E��]������������������������������������������������������������̋�U��j�hP�d�    PQSVW���3�P�E�d�    �e��q������    u�������E�    �Z����$�N����M���   j j ������E������)c��E�����������M�d�    Y_^[��]������������������������������������������������̋�U��Q�E�    �	�E����E��M�U�;}'h���E����M�Q�L�/�������t����2���]���������������������������������̋�U����} t�輿���E��M�}� t�觿���U�:csm�u/�E�xu&�M�y �t�U�z!�t�E�x"�u��h����M�Q�B���E��M�Q�B��M���U����U��E����E��}� ~0�M���U��E��H��Q�M����P��������u�   ��3���]�����������������������������������������������������������U���SQ�E���E��EU�u�M�m������VW��_^��]�MU���   u�   Q����]Y[�� �������������������̋�U������3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ��������UR��������E�P�MQ��������UR��������E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR�0�����f�E�f��f�E��؋Mf�U�f�Q
�M�3�������]����������������������������������������������������������������������������������������������̋�U��=L� uj �EP�MQ�URh��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h��d�    P��H���3�P�E�d�    �EP�M������E�    �} t�M�U�3��} ���Ẽ}� uh��j j^hH�j��������u̃}� uD�����    j j^hH�h4�h���������E�    �E������M��Y����E��  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uhЖj j_hH�j�p�������u̃}� uD�#����    j j_hH�h4�hЖ�&������E�    �E������M�������E��v  �M�M��E�    �U���E�M����M��M��H�����t0�M��<�������   ~�M��)���Pj�E�P�������E��j�M�Q�M�����P�x������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} |�}t�}$~.�} t�U�E��E�    �E������M������E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M����M��U���E�M����M�����3��u�E�j�U�R�M�芼��P���������t�E��0�E��Qh  �M�Q�M��_���P�Ҷ������t0�U��a|�E��z�M�� �M���U�U��E���7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M���U�E����E��!����M����M��U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4������ "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U���E��t�M��ىMЋUЉU��E������M��H����E��M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U��=L� uj�EP�MQ�URh���������j�EP�MQ�URj �n�����]�������������������������̋�U��j�EP�MQ�UR�EP�4�����]���������������̋�U��=L� uj �EP�MQ�URh��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h��d�    P��lVW���3�P�E�d�    �EP�M�������E�    �} t�M�U�3��} ���E��}� uh��j j^h�j�ĸ������u̃}� uN�w����    j j^h�hܗh���z������E�    �E�    �E������M������E��U��<  �} t�}|�}$~	�E�    ��E�   �U��U��}� uhЖj j_h�j�$�������u̃}� uN������    j j_h�hܗhЖ��������E�    �E�    �E������M��p����E��U��  �M�M��E�    �E�    �U���E�M����M��M�������t0�M��߶������   ~�M��̶��Pj�E�P�;������E��j�M�Q�M�訶��P�������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E����E��M���U�E����E��E�RPj�j������E�U�j�M�Q�M�裵��P��������t�U��0�U��Th  �E�P�M��x���P��������t0�M��a|�U��z�E�� �E���M�M��U���7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u^�U�;U�uV�u�3��E�RPj�j������u��}��E��U��E�;E�w.r�M�;M�w$�E�RP�U�R�E�P致���M�3��։EĉU���U���U�} u��E���M�U����U�������E����E��M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI����� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M���U��t�E��؋Mȃ� �ىEĉMȋUĉU��EȉE��E������M�������E��U��M�d�    Y_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�t�����]���������������̋�U��=L� uj�EP�MQ�URh��:�������j�EP�MQ�URj ������]�������������������������̋�U��j�EP�MQ�UR�EP�������]���������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����'  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tE�U�;U�u.�E�H��  ����ًU��  �����;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���(  ���3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T����K���ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �������|���3Ƀ} ����0�����0��� u!h�Dj h  h�Dj��������u̃�0��� uI�����    j h  h�Dh��h�D������ǅ ���������T����:����� �����7  �E��,�����,����Q��@��   ��,���P��������(�����(����t-��(����t$��(�������(��������@��\����
ǅ\���P���\����H$�����х�uV��(����t-��(����t$��(�������(��������@��X����
ǅX���P���X����B$�� ���ȅ�tǅT���    �
ǅT���   ��T�����$�����$��� u!h0Cj h  h�Dj�t�������u̃�$��� uI�$����    j h  h�Dh��h0C�$�����ǅ����������T���������������T6  3Ƀ} ���� ����� ��� u!h�j h  h�Dj��������u̃� ��� uI�����    j h  h�Dh��h�������ǅ����������T����7�����������5  ǅL���    �E������ǅ@���    ���@�������@�����@����q5  ��@���u������ u�Z5  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Uǅ��������ǅ��������ǅp�������ǅ���������E���G�����G����E���E����1  ��L��� ��1  ��G����� |%��G�����x��G�����������P����
ǅP���    ��P�����H�����H���k�	��8�����������8�����8�����  �E���%��  �������u\j
��t���R�EP��������~9��t������$u+��@��� uh@  j ������P袪����ǅ����   �
ǅ����    �������)  j
��t���Q�UR����������������t������E��@��� ��   ������ |#��t������$u������d}ǅL���   �
ǅL���    ��L������������� u!h�j hQ  h�Dj��������u̃���� uI�����    j hQ  h�Dh��h�������ǅ����������T����T�����������2  ������;�x���~��������H������x�����H�����H�����x����   ��8�����   3�tǅD���   �
ǅD���    ��D������������� u!h��j h]  h�Dj��������u̃���� uI������    j h]  h�Dh��h���ο����ǅ����������T����l�����������1  ��8�����@�����@�����.  ��@����$� ���@��� u	������t��@���u�������u�.  ǅ����    ��T���谦��P��G���R�6���������   ��L���P�MQ��G���R�9A  ���E���G����U���U��G�������؉����u!hCj h�  h�Dj��������u̃���� uI�����    j h�  h�Dh��hC蚾����ǅ����������T����8�����������0  ��L���R�EP��G���Q�@  ���-  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �P-  ��G�����<�����<����� ��<�����<���wi��<�����X��$�@����������������D���������������3���������������"�������   ����������������������,  ��G�����*��  ������ u�EP�V������������^  j
��t���Q�UR�ѩ��������������t������E��@��� ��  ������ |#��t������$u������d}ǅ8���   �
ǅ8���    ��8������������� u!h؟j h�  h�Dj���������u̃���� uI�q����    j h�  h�Dh��h؟�q�����ǅ����������T��������������.  ������;�x���~��������4������x�����4�����4�����x����������������� uE��������Ǆ����   ����������G������������������������������   ������P��G���Qj��������������P����������؉����u!h0�j h�  h�Dj芣������u̃���� uI�:����    j h�  h�Dh��h0��:�����ǅ����������T���������������j-  �\*  �+������������������������Q������������������ }���������������������؉������������k�
��G����DЉ�������)  ǅd���    ��)  ��G�����*��  ������ u�UR�r�������d����^  j
��t���P�MQ����������p�����t������U��@��� ��  ��p��� |#��t������$u������d}ǅ0���   �
ǅ0���    ��0������������� u!hx�j h�  h�Dj�ݡ������u̃���� uI�����    j h�  h�Dh��hx�荹����ǅ����������T����+����������+  ��p���;�x���~��p�����,������x�����,�����,�����x�����p����������� uE��p�����Ǆ����   ��p�������G�����������p������������������   ������R��G���Pj��p�����������R� ���������؉� ���u!hНj h�  h�Dj覠������u̃� ��� uI�V����    j h�  h�Dh��hН�V�����ǅ����������T���������������*  �x'  �+��p�����������������������P��������d�����d��� }
ǅd����������d���k�
��G����DЉ�d����'  ��G�����(�����(�����I��(�����(���.�B  ��(��������$�l��U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅ8���    �*����"�������� �������������   �������%  ��G�����$�����$�����A��$�����$���7��"  ��$�������$�����������0  u������   ��������������  �_  ǅ����    ������ u�UR腳����f��<�����  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!hp�j h�  h�Dj臝������u̃����� uI�7����    j h�  h�Dh��hp��7�����ǅ����������T����ս���������g'  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�ѧ��������؉�����u!hȜj h�  h�Dj�w�������u̃����� uI�'����    j h�  h�Dh��hȜ�'�����ǅ����������T����ż���������W&  �   �,��������������������������P荱����f��<�����<���Qh   ��P���R������P�߼���������������� t
ǅl���   �*  ������ u�MQ胸����f��������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hp�j h�  h�Dj�2�������u̃����� uI�����    j h�  h�Dh��hp�������ǅ����������T���耻���������%  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�|���������؉�����u!h(�j h�  h�Dj�"�������u̃����� uI�ҹ���    j h�  h�Dh��h(��ұ����ǅ����������T����p����������$  �j  �,��������������������������R苶����f��������������P���ǅ����   ��P����������  ������ u�UR�H�������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hp�j h�  h�Dj���������u̃����� uI訸���    j h�  h�Dh��hp�訰����ǅ����������T����F�����������"  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�B���������؉�����u!h��j h�  h�Dj��������u̃����� uI蘷���    j h�  h�Dh��h��蘯����ǅ����������T����6�����������!  �0  �+��������������������������P�Q����������������� t�������y u#�`�������������P�k������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������a  ������%0  u��������   ��������d����uǅ���������d������������������������� u�MQ�H�������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hp�j h6  h�Dj���������u̃����� uI訵���    j h6  h�Dh��hp�設����ǅ����������T����F�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�B���������؉�����u!h��j h:  h�Dj��������u̃����� uI蘴���    j h:  h�Dh��h��蘬����ǅ����������T����6�����������  �0  �+��������������������������R�Q�����������������%  tx������ u�d�������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������i������ u�`�����������������������������������������t���������t���������������ɋ�����+������������  ������ u�UR�C�������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hp�j h�  h�Dj��������u̃����� uI裲���    j h�  h�Dh��hp�裪����ǅ����������T����A�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�=���������؉�����u!h��j h�  h�Dj��������u̃����� uI蓱���    j h�  h�Dh��h��蓩����ǅ����������T����1�����������  �+  �+��������������������������P�L������������;�������   3�tǅ���   �
ǅ���    ����������������� u!h�Bj h�  h�Dj��������u̃����� uI貰���    j h�  h�Dh��h�B貨����ǅ����������T����P�����������  �J  �������� t������f��L���f����������L����ǅl���   �  ǅh���   ��G����� ��G�����������@��������������  ��@��� ��  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hp�j h�  h�Dj�Џ������u̃����� uI耯���    j h�  h�Dh��hp�耧����ǅ����������T��������������  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�'���������؉�����u!h��j h�  h�Dj�͎������u̃����� uI�}����    j h�  h�Dh��h���}�����ǅ����������T��������������  �  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��G�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Zh�  htBj��d�����]  R躇���������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�U���U�E�H��P��������������  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!hp�j h  h�Dj�$�������u̃����� uI�Ԭ���    j h  h�Dh��hp��Ԥ����ǅ����������T����r����������  ��@���t!h��j h  h�Dj訌������u̋����������������������������������������H��P���������������T���訋��P��h���P��d���Q��G���R��P���P������Q������R��P��!�Ѓ���������   t-��d��� u$��T����I���P������R��P��!�Ѓ���G�����gu3��������   u%��T�������P������P��Q��!�Ѓ����������-u!��������   ��������������������������P袏������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ��������   t ƅ����0��4�����Q������ǅ����   �*ǅ����   ��������   t��������   ������������% �  �#  ������ u�MQ莓������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u!hp�j h�  h�Dj��������u̃�l��� uI�ʩ���    j h�  h�Dh��hp��ʡ����ǅ����������T����h�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�d���������؉�h���u!h��j h�  h�Dj�
�������u̃�h��� uI躨���    j h�  h�Dh��h��躠����ǅ����������T����X�����������  �R  �1����������������d�����d���R葑������x�����|�����
  ������%   �#  ������ u�MQ�Z�������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������`�����`��� u!hp�j h�  h�Dj��������u̃�`��� uI薧���    j h�  h�Dh��hp�薟����ǅ����������T����4�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�0���������؉�\���u!hH�j h�  h�Dj�ֆ������u̃�\��� uI膦���    j h�  h�Dh��hH�膞����ǅ����������T����$����������  �  �1����������������X�����X���R�]�������x�����|�����  �������� �a  ��������@�'  ������ u�UR�����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������T�����T��� u!hp�j h�  h�Dj装������u̃�T��� uI�S����    j h�  h�Dh��hp��S�����ǅ����������T��������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�P���u!h(�j h�  h�Dj蓄������u̃�P��� uI�C����    j h�  h�Dh��h(��C�����ǅ����������T��������������s  ��  �3����������������L�����L���P�����������x�����|����&  ������ u!�MQ�Ԡ���������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������H�����H��� u!hp�j h�  h�Dj�z�������u̃�H��� uI�*����    j h�  h�Dh��hp��*�����ǅ����������T����ȣ���������Z  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�č��������؉�D���u!h(�j h�  h�Dj�j�������u̃�D��� uI�����    j h�  h�Dh��h(�������ǅ����������T���踢���������J  �  �5����������������@�����@���R�Ӟ���������x�����|����V  ��������@�%  ������ u�MQ蚞�������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������<�����<��� u!hp�j h  h�Dj�C�������u̃�<��� uI�����    j h  h�Dh��hp�������ǅ����������T���葡���������#  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q荋��������؉�8���u!h(�j h  h�Dj�3�������u̃�8��� uI�����    j h  h�Dh��h(�������ǅ|���������T���聠����|����
  �{  �2����������������4�����4���R蜜�������x�����|����"  ������ u�EP�u�����3ɉ�x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������0�����0��� u!hp�j h0  h�Dj�������u̃�0��� uI�͞���    j h0  h�Dh��hp��͖����ǅx���������T����k�����x�����  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�g���������؉�,���u!h(�j h4  h�Dj�~������u̃�,��� uI轝���    j h4  h�Dh��h(�轕����ǅt���������T����[�����t�����  �U  �3����������������(�����(���R�v�����3ɉ�x�����|�����������@tG��|��� >|	��x��� s3��x����؋�|����� �ى�p�����t�����������   ���������x�����p�����|�����t����������� �  u(������%   u��p�����t����� ��p�����t�����d��� }ǅd���   �%�����������������d���   ~
ǅd���   ��p����t���u
ǅ����    ��O�����������d�����d�������d�������p����t�����   �������RP��t���P��p���Q�E�����0�������������RP��t���R��p���P�T�����p�����t���������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�s  ��l��� �B  ��������@t[��������   tƅ����-ǅ����   �:��������tƅ����+ǅ����   ���������tƅ���� ǅ����   ������+�����+�������$�����������u��L���Q�UR��$���Pj �m  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��$���Qj0�  �������� ��   ������ ��   ǅ���    �������� �����������������������������������   �� ���f�f������������Rj�����P�����Q�Ś����������� ������� �������� u	����� uǅL��������-��|���P��L���Q�UR�����P�����Q�  ���S����(��|���R��L���P�MQ������R������P�P  ����L��� |'��������t��L���R�EP��$���Qj ��  �������� tj������R�;�����ǅ����    ������8��� t��8���tǅ����    �
ǅ����   ���������������� u!hؘj h�  h�Dj�tx������u̃���� uI�$����    j h�  h�Dh��hؘ�$�����ǅp���������T��������p����T  �������%  ��@��� �  ǅ����    ���������������������;�x�����  �����������������������������������������  �������$�$����������E�������MQ�d������  ���������E�������MQ�������_  ���������E�������MQ�������;  ���������E�������MQ�������  ���������E�������MQ��������   ���������E�������MQ谓������   ���������E�������MQ�z������h�����l����   3�tǅ����   �
ǅ����    ���������������� u!hh�j h.	  h�Dj�Dv������u̃���� uF������    j h.	  h�Dh��hh�������ǅd���������T���蒖����d����'������s�����L�����`�����T����i�����`����M�3�������]Ë�8�f���J��.���`��#����6�E� �I i�9�-�J�[� �m������h�����~�m����;�����}�   	
B�f�����Ұ��J���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�}�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U���<  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��0q���E�    �+����E�3Ƀ} �������������� u!h�Dj h  h�Dj�1c������u̃����� uF�����    j h  h�Dh$�h�D��z����ǅ��������M�肃��������#  �E�������������Q��@��   ������P�do�����������������t-�������t$�������������������@�������
ǅ����P��������H$�����х�uV�������t-�������t$�������������������@�������
ǅ����P��������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h0Cj h  h�Dj�a������u̃����� uF�l����    j h  h�Dh$�h0C�ly����ǅ��������M�����������  3Ƀ} �������������� u!h�j h  h�Dj�4a������u̃����� uF�����    j h  h�Dh$�h���x����ǅ��������M�腁��������&  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���  ������ �	  �������� |%��������x�������������������
ǅ����    ������������������k�	��������������������������   3�tǅ����   �
ǅ����    ������������������ u!h��j ha  h�Dj��_������u̃����� uF�x���    j ha  h�Dh$�h���xw����ǅ��������M�����������  ��������������������  �������$�0��E�    �M��^��P������R�a��������   ������P�MQ������R�u  ���E��������U���U����������؉�|���u!hCj h�  h�Dj��^������u̃�|��� uF�v~���    j h�  h�Dh$�hC�vv����ǅ��������M����������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK��������h��$�P��E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�~z�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�%z�����Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  �����������$�|��E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  �����������$����U���0  u�E�   �E��M���  tUǅx���    �UR��p����f������������Ph   ������Q�U�R�M|������x�����x��� t�E�   �&�EP� x����f��t�����t����������E�   �������U��W  �EP��w������p�����p��� t��p����y u�`��U��E�P��^�����E��P�M���   t&��p����B�E���p�����+����E��E�   ��E�    ��p����B�E���p�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������h����MQ��v�����E��U���  te�}� u�d��E��E�   �M���d�����h�����h�������h�����t��d������t��d�������d����ɋ�d���+M����M��[�}� u	�`��U��E���l�����h�����h�������h�����t��l������t��l�������l����ɋ�l���+E��E��  �MQ�v������`����	j������   3�tǅ����   �
ǅ����    ��������\�����\��� u!h�Bj h�  h�Dj��X������u̃�\��� uF�x���    j h�  h�Dh$�h�B�p����ǅ ��������M��!y���� �����  ��  �U��� t��`���f������f����`�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  htBj�Ú�]  R�Q�����E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���P�����T����M��V��P�E�P�M�Q������R�E�P�M�Q��P���R��P��!�Ѓ��M���   t$�}� u�M��kV��P�U�R��P��!�Ѓ���������gu*�U���   u�M��6V��P�E�P��Q��!�Ѓ��U����-u�M���   �M��U����U��E�P��Z�����E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�_������@�����D����   �U���   t�EP��^������@�����D����   �M��� tB�U���@t�EP�r��������@�����D�����MQ�r���������@�����D����=�U���@t�EP�\r�������@�����D�����MQ�Ar����3҉�@�����D����E���@t@��D��� 7|	��@��� s,��@����ً�D����� �ډ�8�����<����E�   �E����@�����8�����D�����<����E�% �  u&�M���   u��8�����<����� ��8�����<����}� }	�E�   ��M�����M��}�   ~�E�   ��8����<���u�E�    �E��E��M̋Ũ��U̅���8����<���t{�E��RP��<���Q��8���R�Kt����0��L����E��RP��<���P��8���Q�]r����8�����<�����L���9~��L����������L����E���L�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅4����M���u������R�EP��4���Qj �K	  ���U�R������P�MQ�U�R�E�P�|	  ���M���t$�U���u������P�MQ��4���Rj0� 	  ���}� ��   �}� ��   ǅ���    �E���0����M܉�,�����,�����,�������,�������   ��0���f�f������������Pj�� ���Q��(���R�^s�����������0�������0�������� u	��(��� uǅ���������*�M�Q������R�EP��(���Q�� ���R�{  ���V�����E�P������Q�UR�E�P�M�Q�U  �������� |$�U���t������P�MQ��4���Rj ��  ���}� tj�E�P��d�����E�    ����������� t������tǅ����    �
ǅ����   ���������������� u!hؘj h�  h�Dj�%Q������u̃���� uC��p���    j h�  h�Dh$�hؘ��h����ǅ���������M��vq����������������������M��Zq���������M�3��t����]ÍI ������/�|������	������!�*� �I 7������� ���C���]�����Y�;�����V���M�i�D�   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�]b�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    �E������E�    j�C������u����C  j��I�����E�    �E�    �	�E���E�}�@��  �M�<�@ �#  �U��@�E��	�M؃�@�M؋U��@   9E���   �M��Q����   �E؃x uaj
�_I�����E�   �M؃y u.h�  �U؃�R�D"��u	�E�   ��E؋H���U؉J�E�    �   �j
��Y����Ã}� u+�E؃�P��"�M��Q��t�E؃�P��"�4����}� u-�M��A�U�������E����M�U�+�@��E��������}��t��   ��   h�   h@�jj@j �e�����E؃}� ��   �E�M؉�@���� ���	�E؃�@�E؋M��@��   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃�����@�D�U�R��A������u�E������������E������   �j�X����ËE܋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} ��   �E;���   �M���U������@�<�um�=�uB�M�M��}� t�}�t�}�t�(�URj��#��EPj��#��MQj��#�U���E������@�U�3����Od��� 	   �jM���     �����]�����������������������������������������������������������̋�U��Q�} ��   �E;���   �M���U������@�L����   �U���E������@�<�th�=�u<�U�U��}� t�}�t�}�t�"j j��#�j j��#�
j j��#�E���M������@�����3����0c��� 	   �KL���     �����]������������������������������������������������������������̋�U����}�u��K���     �b��� 	   ����2  �} |�E;�s	�E�   ��E�    �M�M��}� u!h@~j h;  h��j�B������u̃}� u<�}K���     �Lb��� 	   j h;  h��h|�h@~�LZ��������   �E���M������@�D
������؉E�u!h|}j h<  h��j�B������u̃}� u9��J���     ��a��� 	   j h<  h��h|�h|}��Y���������U���E������@���]����������������������������������������������������������������������������������������������̋�U��j�h@�h)d�    P���SVW���1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP�H"�E��}� u�$"P�,>��������q  �}�u�M��@�M���}�u
�U���U��vb���E؃}��u�B`���    �]I���     ����#  �E�    �EP�M�Q�*d�����U���U�E����M؃�����@�E�D
�M����U؃�����@�L$�ဋU����E؃�����@�L$�E����M؃�����@�D
$$�M����U؃�����@�D$�E�   �E������   �K�}� u8�U����E؃�����@�T����E����M؃�����@�T�M�Q� ;����Ã}� t�U؉U���E������EԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h`�h)d�    P���SVW���1E�3�P�E�d�    �E���M�����@�M��E�   �U��z u_j
��?�����E�    �E��x u,h�  �M���Q�D"��u�E�    �U��B���M��A�E������   �j
�|P����Ã}� t!�U���E������@�TR��"�E�M�d�    Y_^[��]��������������������������������������������������������������������������̋�U��E���M������@�D
P��"]������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    j�>�����E�    �EP�5\����f�E��E������   �j�IO�����f�E�M�d�    Y_^[��]���������������������������������������������̋�U��Q�=���u�V7���=���u���  �(j �E�Pj�MQ���R��"��u���  �f�E��]��������������������������������̋�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M��oI���M���:������   t1�M���:��� ���   th��j jGh�j�t;������u̍M��:����z u*�} t�Ef��Uf�
�E�   �M���[���E��R  �M��z:��P�E�Q�=��������   �M��Z:������   ~R�M��G:��� �M;��   |=3҃} ��R�EP�M��$:������   R�EPj	�M��:����QR��!��uB�M���9��� �M;��   r�U�B��u"�NZ��� *   �E������M��[���E��   �M��9������   �U�M���Z���E��k�a3��} ��P�MQj�URj	�M��{9��� �HQ��!��u��Y��� *   �E������M��Z���E���E�   �M��Z���E���M��}Z����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR��V����]�������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�    j�:�����E�    �E�   �	�E����E��M�;���   �U�l��<� t|�M��l����H��   t"�U�l���Q�7�������t	�U���U�}�|=�E��l����� R�P"j�E��l���R�K�����E��l���    �Y����E������   �j�J����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �} uj �  ���@�EP��F�����E�    �MQ��N�����E��E������   ��UR�M����ËE�M�d�    Y_^[��]������������������������������������������̋�U��} uj �n  ���@�EP�S������t����+�M�Q�� @  t�EP�TC����P�&@��������3�]�����������������������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R��B����P�5����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����������������������������������������������������̋�U��j�   ��]���������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j��6�����E�    �E�    �	�E����E��M�;���   �U�l��<� ��   �M��l����H��   ��   �U�l���Q�U�R�W�����E�   �E��l����B%�   te�}u%�M��l���P�L�������t	�M���M��:�} u4�U�l����Q��t!�E��l���R��K�������u�E������E�    �   ��E��l���R�E�P�J�����������E������   �j�F����Ã}u�E����E܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������̋�U����} uh�Aj j?hȤj�23������u̋M�M��U�R��?����P��K������u3��  �.D���� 9E�u	�E�    ��D����@9E�u	�E�   �3���   �X����X��M��Q��  t3��   �E��<�`� u\j[h��jh   �g,�����E�M��U��`��}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U���`��A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]��������������������������������������������������������������������������������������̋�U��Q�} t'�}t!h@�j h�   hȤj�{1������u̋M�M��} tG�U��B%   t:�M�Q�8N�����U��B%�����M��A�U��B    �E��     �M��A    ��]��������������������������������������̋�U��j�h�h)d�    P���SVW���1E�3�P�E�d�    ��A���� �E�3��} ���E؃}� uh�j j4h��j�0������u̃}� u+�DP���    j j4h��hx�h��GH��������i�U�R�?�����E�    �E�P�/�����E܋MQ�UR�EP�M�Q�U���E��U�R�E�P�L�����E������   ��M�Q�kF����ËE��M�d�    Y_^[��]�����������������������������������������������������������������������̋�U��EP�MQ�URhA9�i,����]����������������̋�U��EP�MQ�URh<�9,����]����������������̋�U��EP�MQ�URh=�	,����]����������������̋�U��EPj �MQhA9��+����]������������������̋�U��EPj �MQh<�+����]������������������̋�U��EPj �MQh=�{+����]������������������̋�U���   ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���;���E�    ��M���E�3Ƀ} �������������� u!h�Dj h  h�Dj��-������u̃����� uF�M���    j h  h�Dh�h�D�E����ǅ8��������M��2N����8����  3��} �������������� u!h�j h  h�Dj�Y-������u̃����� uF�	M���    j h  h�Dh�h��	E����ǅ4��������M��M����4����z  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���h  ������ �[  �������� |%��������x�������������� ����
ǅ ���    �� ���������������k�	��������������������������   3�tǅ���   �
ǅ���    ����������������� u!h��j ha  h�Dj��+������u̃����� uF�K���    j ha  h�Dh�h���C����ǅ0��������M��<L����0����  �����������������*  ������$�\
�E�   ������Q�UR������P�Y  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ������������������ ����������wL��������
�$�|
�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�uG�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�G�����Ẽ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  ��������
�$��
�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  �������(�$��
�M���0  u	�U��� �U��E�   �EP�RE����f�������M��� tW���������   ������ƅ���� �M��'��P�M��y'��� ���   Q������R������P��E������}�E�   �f������f�������������U��E�   �  �EP�D���������������� t�������y u�`��U��E�P��+�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ�����������|����MQ��C�����E��U��� ��   �}� u�`��E��M��������E�    �	�U܃��U܋E�;�|���}L���������t?�M���%��P�������Q�z(������t������������������������������d�}� u	�d��M��E�   �U���x�����|�����|�������|�����t��x������t��x�������x����ɋ�x���+U����U��  �EP��B������t�����6������   3�tǅ���   �
ǅ���    �������p�����p��� u!h�Bj h�  h�Dj�%������u̃�p��� uF�ME���    j h�  h�Dh�h�B�M=����ǅ,��������M���E����,����  ��  �M��� t��t���f������f����t�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  htBj�Ḿ�]  Q�V�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��#��P�U�R�E�P������Q�U�R�E�P��h���Q��R��!�Ѓ��E�%�   t%�}� u�M��8#��P�M�Q��R��!�Ѓ���������gu)�M���   u�M��#��P�U�R��P��!�Ѓ��M����-u�E�   �E��M����M��U�R�'�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ��+������X�����\����   �U���   t�EP�+������X�����\����   �M��� tB�U���@t�EP�f?��������X�����\�����MQ�J?���������X�����\����=�U���@t�EP�$?�������X�����\�����MQ�	?����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R�A����0��d����E��RP��T���P��P���Q�"?����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �N  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M����P�M��v������   R��H���P������Q��<������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�v  �������� |$�U���t������P�MQ��L���Rj ��  ���}� tj�E�P�1�����E�    �s��������� t������tǅ ���    �
ǅ ���   �� �����<�����<��� u!hؘj h�  h�Dj��������u̃�<��� uC�=���    j h�  h�Dh�hؘ�5����ǅ(��������M��G>����(������������$����M��+>����$����M�3���@����]�h�����8�������������*�3� �I A������
� ��L�� ����`�m���� ��   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�)0�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����#  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tA�U�;U�u*�E�H�� ��Ƀ��U�� ��҃�;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ���3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T���� ��ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �)2����|���3Ƀ} ����0�����0��� u!h�Dj h  h�Dj�,������u̃�0��� uI��1���    j h  h�Dh8�h�D��)����ǅ,���������T����z2����,����3  3��} ����,�����,��� u!h�j h  h�Dj�������u̃�,��� uI�Q1���    j h  h�Dh8�h��Q)����ǅ(���������T�����1����(����3  ǅL���    �U������ǅ@���    ���@�������@�����@�����2  ��@���u������ u�2  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Mǅ��������ǅ��������ǅp�������ǅ���������Uf�f��D�����D����U���U���K/  ��L��� �>/  ��D����� |%��D�����x��D����������������
ǅ����    ��������H�����H���k�	��8�����������8�����8�����  �U���%��  �������u\j
��t���Q�UR�M������~9��t������$u+��@��� uh@  j ������R�X����ǅ����   �
ǅ����    �������)  j
��t���P�MQ����������������t������U��@��� ��   ������ |#��t������$u������d}ǅ����   �
ǅ����    ��������(�����(��� u!h�j hQ  h�Dj�������u̃�(��� uI�l.���    j hQ  h�Dh8�h��l&����ǅ$���������T����
/����$����40  ������;�x���~���������������x�����������������x����   ��8�����   3�tǅ����   �
ǅ����    ��������$�����$��� u!h��j h]  h�Dj��������u̃�$��� uI�-���    j h]  h�Dh8�h���%����ǅ ���������T����".���� ����L/  ��8����������������N,  �������$��I��@��� u	������t��@���u�������u�,  ǅ����   ��L���Q�UR��D���P�=  ����+  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �+  ��D����������������� ������������wj���������I�$��I���������������E���������������4���������������#�������ʀ   ����������������������	+  ��D�����*��  ������ u�UR��(�����������`  j
��t���P�MQ�y��������������t������U��@��� ��  ������ |#��t������$u������d}ǅ|���   �
ǅ|���    ��|����� ����� ��� u!h؟j h�  h�Dj�Q������u̃� ��� uI�+���    j h�  h�Dh8�h؟�#����ǅ���������T����+���������,  ������;�x���~��������x������x�����x�����x�����x����������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R���������؉����u!h0�j h�  h�Dj�
������u̃���� uI��)���    j h�  h�Dh8�h0���!����ǅ���������T����f*��������+  �(  �+������������������������P�&���������������� }���������������������ډ������������k�
��D����TЉ������2(  ǅd���    �#(  ��D�����*��  ������ u�MQ� &������d����`  j
��t���R�EP���������p�����t������M��@��� ��  ��p��� |#��t������$u������d}ǅt���   �
ǅt���    ��t������������� u!hx�j h�  h�Dj�k������u̃���� uI�(���    j h�  h�Dh8�hx�� ����ǅ���������T����(���������)  ��p���;�x���~��p�����p������x�����p�����p�����x�����p����������� uG��p�����Ǆ����   ��p�����f��D���f��������p������������������   ������Q��D���Rj��p�����������Q���������؉����u!hНj h�  h�Dj�2������u̃���� uI��&���    j h�  h�Dh8�hН������ǅ���������T����'��������(  ��%  �+��p���������������������R�#������d�����d��� }
ǅd����������d���k�
��D����TЉ�d����_%  ��D�����l�����l�����I��l�����l���.�D  ��l�����J�$�J�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������d�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu������   �������ǅ8���    ������#�������� ���������������   ��������#  ��D�����h�����h�����A��h�����h���7�B!  ��h������J�$�HJ��������0  u�������� ������ǅ����   ������ u�EP�v!����f��<�����  ������ |������d}ǅd���   �
ǅd���    ��d������������� u!hp�j hv  h�Dj�%������u̃���� uI��#���    j hv  h�Dh8�hp�������ǅ���������T����s$��������%  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P���������؉����u!h(�j hz  h�Dj�������u̃���� uI��"���    j hz  h�Dh8�h(�������ǅ���������T����a#��������$  �  �,���������������� ����� ���Q�|����f��<����������� t_��<���%�   ������ƅ���� ��T������P��T����������   R������P��P���Q��������}
ǅl���   �f��<���f��P�����P���������ǅ����   �^  ������ u�MQ��������������  ������ |������d}ǅ`���   �
ǅ`���    ��`��������������� u!hp�j h�  h�Dj�}������u̃����� uI�-!���    j h�  h�Dh8�hp��-����ǅ���������T�����!���������"  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q����������؉�����u!h��j h�  h�Dj�k ������u̃����� uI� ���    j h�  h�Dh8�h�������ǅ ���������T���� ���� �����!  �w  �+��������������������������R������������������ t�������x u#�`�������������R�������������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q��������������������  ��������0  u�������� ��������d����uǅ\���������d�����\�����\��������������� u�EP��������������  ������ |������d}ǅX���   �
ǅX���    ��X��������������� u!hp�j h6  h�Dj�~�������u̃����� uI�.���    j h6  h�Dh8�hp��.����ǅ����������T���������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P��	��������؉�����u!h��j h:  h�Dj�l�������u̃����� uI����    j h:  h�Dh8�h�������ǅ����������T��������������  �x  �+��������������������������Q�������������������� ��   ������ u�`�������������������ǅ����    ���������������������;�����}O���������tB��T��������P�������Q�D�������t������������������������������v������ u�d�������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������'  ������ u�EP�������������  ������ |������d}ǅT���   �
ǅT���    ��T��������������� u!hp�j h�  h�Dj�F�������u̃����� uI�����    j h�  h�Dh8�hp�������ǅ����������T�������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P���������؉�����u!h��j h�  h�Dj�4�������u̃����� uI�����    j h�  h�Dh8�h��������ǅ����������T�������������  �@  �+��������������������������Q������������
������   3�tǅP���   �
ǅP���    ��P��������������� u!h�Bj h�  h�Dj�S�������u̃����� uI����    j h�  h�Dh8�h�B�����ǅ����������T��������������  �_  �������� t������f��L���f����������L����ǅl���   �%  ǅh���   ��D����� f��D�����������@��������������  ��@��� ��  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u!hp�j h�  h�Dj� �������u̃����� uI�����    j h�  h�Dh8�hp�������ǅ����������T����n���������  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R���������؉�����u!h��j h�  h�Dj��������u̃����� uI�����    j h�  h�Dh8�h��������ǅ����������T����i���������  �'  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��D�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Yh�  htBj��d���]  P�	����������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�E���E�M�Q��A��������������  ������ |������d}ǅH���   �
ǅH���    ��H��������������� u!hp�j h  h�Dj�s�������u̃����� uI�#���    j h  h�Dh8�hp��#����ǅ����������T���������������  ��@���t!h��j h  h�Dj���������u̋����������������������������������������Q��A���������������T��������P��h���Q��d���R��D���P��P���Q������R������P��Q��!�Ѓ���������   t.��d��� u%��T�������P������P��Q��!�Ѓ���D�����gu2������%�   u%��T����Y���P������Q��R��!�Ѓ����������-u!��������   ��������������������������Q��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ������%�   t&�0   f��������4�����Qf������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  �%  ������ u�EP���������������������  ������ |������d}ǅD���   �
ǅD���    ��D��������������� u!hp�j h�  h�Dj�c�������u̃����� uI����    j h�  h�Dh8�hp��
����ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�����������؉�����u!h��j h�  h�Dj�Q�������u̃����� uI����    j h�  h�Dh8�h���	����ǅ����������T��������������  �]  �1��������������������������Q��������������������  ��������   �%  ������ u�EP��������������������  ������ |������d}ǅ@���   �
ǅ@���    ��@��������������� u!hp�j h�  h�Dj�,�������u̃����� uI�����    j h�  h�Dh8�hp�������ǅ����������T����z���������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P����������؉�|���u!hH�j h�  h�Dj��������u̃�|��� uI�����    j h�  h�Dh8�hH�������ǅ����������T����h���������  �&  �1����������������x�����x���Q��������������������  �������� �e  ��������@�)  ������ u�MQ�?��������������������  ������ |������d}ǅ<���   �
ǅ<���    ��<�����t�����t��� u!hp�j h�  h�Dj���������u̃�t��� uI����    j h�  h�Dh8�hp������ǅ����������T����5���������_  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�V���������؉�p���u!h(�j h�  h�Dj���������u̃�p��� uI����    j h�  h�Dh8�h(������ǅ����������T����#���������M  ��  �3����������������l�����l���R�>	�������������������(  ������ u!�EP�	���������������������  ������ |������d}ǅ8���   �
ǅ8���    ��8�����h�����h��� u!hp�j h�  h�Dj��������u̃�h��� uI�l���    j h�  h�Dh8�hp��l����ǅ����������T����
���������4  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�+���������؉�d���u!h(�j h�  h�Dj��������u̃�d��� uI�Z
���    j h�  h�Dh8�h(��Z����ǅ����������T�����
���������"  �  �5����������������`�����`���Q���������������������Z  ��������@�'  ������ u�EP���������������������  ������ |������d}ǅ4���   �
ǅ4���    ��4�����\�����\��� u!hp�j h  h�Dj��������u̃�\��� uI�3	���    j h  h�Dh8�hp��3����ǅ����������T�����	����������
  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�����������؉�X���u!h(�j h  h�Dj�q�������u̃�X��� uI�!���    j h  h�Dh8�h(��! ����ǅ����������T��������������	  �}  �2����������������T�����T���Q��������������������$  ������ u�UR�����3ɉ�������������  ������ |������d}ǅ0���   �
ǅ0���    ��0�����P�����P��� u!hp�j h0  h�Dj�[�������u̃�P��� uI����    j h0  h�Dh8�hp�������ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�����������؉�L���u!h(�j h4  h�Dj�I�������u̃�L��� uI�����    j h4  h�Dh8�h(��������ǅ����������T��������������  �U  �3����������������H�����H���R�����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ��������������d��� }ǅd���   �%�����������������d���   ~
ǅd���   �����������u
ǅ����    ��O�����������d�����d�������d������������������   �������RP������P������Q�����0�������������RP������R������P���������������������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�k  ��l��� �:  ��������@tj��������   t�-   f������ǅ����   �D��������t�+   f������ǅ����   �!��������t�    f������ǅ����   ������+�����+�������D�����������u��L���Q�UR��D���Pj ��  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��D���Qj0�  �������� ��   ������ ��   ��������@�����������<�����<�����<�������<�������   ��T����Y���P��T����M���� ���   Q��@���R��<���P��������8�����8��� ǅL��������2��L���Q�UR��<���P�E  ����@����8�����@����`����(��|���R��L���P�MQ������R������P��  ����L��� |'��������t��L���R�EP��D���Qj �T  �������� tj������R������ǅ����    ������8��� t��8���tǅ,���    �
ǅ,���   ��,�����4�����4��� u!hؘj h�  h�Dj��������u̃�4��� uI�h ���    j h�  h�Dh8�hؘ�h�����ǅ����������T�������������0  �������  ��@��� ��  ǅ����    ���������������������;�x�����  ����������������(�����(�������(�����(�����   ��(����$��J���������E�������MQ�������_  ���������E�������MQ�������;  ���������E�������MQ�~������  ���������E�������MQ�Z�������   ���������E�������MQ��������   ���������E�������MQ�������������������   3�tǅ$���   �
ǅ$���    ��$�����0�����0��� u!hh�j h.	  h�Dj��������u̃�0��� uF�\����    j h.	  h�Dh8�hh��\�����ǅ����������T���������������'�����#�����L�����������T���������������M�3������]Ë���&���d!�"��p_�� �I �!�"�!�"�" �/#�(g4�%7/0#04,�4]4�(N4s4AD   	
�G"HFHjH�H�H�H�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U��j�h0�h)d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� uhܦj j3hh�j�\�������u̃}� u-�����    j j3hh�hX�hܦ���������  �M�U�U�E�P�z������E�    �M�Q�UR�c�����f�E��E������   ��E�P�Q������f�E��M�d�    Y_^[��]����������������������������������������������������������������������������̋�U���8���3ŉE�V�E�H��@�d  �UR����������t@�EP����������t/�MQ������������UR������������@�E���E�P��E�H$�����у�tj�EP���������t@�MQ���������t/�UR�p����������EP�_����������@�E���E�P��M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ�D������  �(  �UR����������t@�EP���������t/�MQ�����������UR�����������@�E���E�P��E��H��   ��   �URj�E�P�M�Q��������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R�T������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP������^�M�3��������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�D�����]��������̋�U���8�EP�M��Q���3Ƀ} ���M�}� uh�\j j4h �j�j�������u̃}� u=�����    j j4h �h �h�\� ������E�����M�������E��  3��} ���E��}� uh�[j j5h �j���������u̃}� u=�����    j j5h �h �h�[�������E�����M��Q����E��   �M��������z u"�EP�MQ��������EԍM������E��x�b�U��E̍M�����P�M�Q�V������E��U���U�E��MȍM�����P�U�R�,������E��E���E�}� t�M�;M�t��U�+U��UЍM������EЋ�]����������������������������������������������������������������������������������������������������������̋�U����E��M��U��E���E��A|�}�Z	�M��� �M��U��E��M��U���U��A|�}�Z	�E��� �E��}� t�M�;M�t��E�+E���]������������������������������̋�U����=L� ��   3��} ���E��}� uh�\j jbh �j���������u̃}� u0�|����    j jbh �h��h�\�����������   3҃} �U��}� uh�[j jch �j�c�������u̃}� u-�����    j jch �h��h�[�����������&�MQ�UR�h�������j �EP�MQ��������]������������������������������������������������������������������������̋�U���@�} �!  �EP�M��W���3Ƀ} ���M�}� uh�\j j;h��j�p�������u̃}� u=�#����    j j;h��hاh�\�&������E�����M�������E��  3��} ���E��}� uh�[j j<h��j���������u̃}� u=�����    j j<h��hاh�[�������E�����M��W����E��1  ����;U����E�uh��j j=h��j��������u̃}� u=�=����    j j=h��hاh���@������E�����M�������E��   �M�������z u)�EP�MQ�UR�7������E̍M������E��   �m�E��MčM��E���P�U�R��������E��E���E�M��U��M�����P�E�P�������E��M���M�U���Ut�}� t�E�;E�t��M�+M��MȍM��%����E��3���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����=L� �Y  3��} ���E��}� u!h�\j h�   h��j��������u̃}� u3�Y����    j h�   h��hp�h�\�Y����������  3҃} �U��}� u!h�[j h�   h��j�:�������u̃}� u3������    j h�   h��hp�h�[������������   ����;M҃��U�u!h��j h�   h��j���������u̃}� u0�����    j h�   h��hp�h�������������.�MQ�UR�EP蘺������j �MQ�UR�EP��������]��������������������������������������������������������������������������������������������������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   ����}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q��!_^��]� ���������������������̋�U��Q�M��E�� ���M��A    �U��B �E���]����������������������̋�U��Q�M��M��j����E��t�M�Q��������E���]� �����������������̋�U��Q�M��E�� ���M��A    �U��B �E�Q�M�艺���E���]� ���������������������̋�U��Q�M��E�� ���M��U��A�M��A �E���]� ������������������̋�U��Q�M��E�� ���M��A    �U��B �EP�M�������E���]� �����������������������̋�U��Q�M��E�;Et0�M�諻���M�Q��t�E�HQ�M�觹����U��E�H�J�E���]� ���������������������̋�U��Q�M��E�� ���M��J�����]������������������̋�U����M��E��x t�M��Q�U���E����E���]�������������������̋�U����M��} tK�EP����������E��M�Q��������U��B�E��x t�MQ�U�R�E��HQ�������U��B��]� �����������������������������̋�U��Q�M��E��H��t�U��BP��������M��A    �U��B ��]������������������������̋�U��Q�M��EP�M��r����M��ܨ�E���]� ��������̋�U��Q�M��M������E��t�M�Q�ӽ�����E���]� �����������������̋�U��Q�M��EP�M��!����M��ܨ�E���]� ��������̋�U��Q�M��E�� ܨ�M�������]������������������̋�U��Q�M��EP�M������M����E���]� ��������̋�U��Q�M��M��V����E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M��Q����M����E���]� ��������̋�U��Q�M��E�� ��M��1�����]������������������̋�U��Q�M��EP�M��z����M�����E���]� ��������̋�U��Q�M��M�������E��t�M�Q�3������E���]� �����������������̋�U��Q�M��EP�M��E����M�����E���]� ��������̋�U��Q�M��E�� ���M�������]������������������̋�U��j j jj jh   @h��#���]����������̋�U��=���t�=���t���P�#]�����������̋�U��j�hP�h)d�    P���SVW���1E�3�P�E�d�    �E�����3��} ���E��}� uh�Dj j.h0�j�Ÿ������u̃}� u+�x����    j j.h0�h�h�D�{���������W�U�B��@t�M�A    �=�UR��������E�    �EP�:������E��E������   ��MQ������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U����E�����3��} ���E�}� uhܦj jYh0�j蟷������u̃}� u.�R����    j jYh0�h��hܦ�U���������   �U�U��E��H��   ta�U�R�-������E��E�P臻�����M�Q�������P��������}	�E������$�U��z tj�E��HQ�Z������U��B    �E��@    �E���]�����������������������������������������������������������������������̋�U��j�hp�h)d�    P���SVW���1E�3�P�E�d�    �}�u����� 	   ����  �} |�E;�s	�E�   ��E�    �M؉M��}� uh��j j,h �j��������u̃}� u.����� 	   j j,h �h�h������������;  �E���M������@�D
������؉E�uhȩj j-h �j荵������u̃}� u.�@���� 	   j j-h �h�hȩ�C����������   �UR�������E�    �E���M������@�D
��t;�MQ�������P�#��u�$"�E���E�    �}� u�>�Խ���U������ 	   �E�����3�uh�|j jEh �j跴������u��E������   ��UR�<�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�   ��]�������������������̋�U���$�} t�E�M�3҃} �U�}� uh��j j^h8�j舳������u̃}� u-�;����    j j^h8�h �h���>�����3��'  �} t�}|�}$~	�E�    ��E�   �M��M�}� uhЖj j_h8�j�	�������u̃}� u-�����    j j_h8�h �hЖ������3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q�3�������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R��������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q�կ������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q臯�����E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4�<���� "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�X�����]�������������������̋�U��j�EP�MQ�UR�(�����]�������������������̋�U��j�EP�MQ�UR�������]�������������������̋�U��� �} uh�Aj jdhXAj肮������u̋M�M��U�R�������E��E��H��   u&����� 	   �U��B�� �M��A���  �c  �/�U��B��@t$������ "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6蕾���� 9E�t舾����@9E�u�M�Q�)�������u�U�R�j������E��H��  �  �U��E��
+Hy!h�@j h�   hXAj���������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�#������E��s�}��t!�}��t�M����U������@�U���E�P��E��H�� t9jj j �U�R�6������E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q�o������E�U�;U�t�E��H�� �U��J���  ��E%��  ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̋�U��j�h��h)d�    P���SVW���1E�3�P�E�d�    �}�u�E����     ����� 	   ����  �} |�E;�s	�E�   ��E�    �M؉M��}� uh@~j j.h��j���������u̃}� u9�ֲ���     ����� 	   j j.h��h��h@~����������  �E���M������@�D
������؉E�uh|}j j/h��j�w�������u̃}� u9�P����     ����� 	   j j/h��h��h|}�"���������   �UR�Ƥ�����E�    �E���M������@�D
��t�MQ�H������E��4����� 	   �E�����3�uh�|j j9h��j���������u��E������   ��MQ�E�����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QV�EP辵�������t]�}u�@���   ��u�}u(�@�HD��tj胵������j�w�����;�t�UR�g�����P�#��t	�E�    �	�$"�E��EP�������M���U������@�D �}� t�M�Q詤��������3�^��]����������������������������������������������������̋�U��} uh��j j.h0�j�զ������u̋M�Q��   tK�E�H��t@j�U�BP�������M�Q�������E�P�M�    �U�B    �E�@    ]��������������������������������������������̋�U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%�!�%�!�%�!�%�!�%�!�%�!�%�!�%�!�%�!�%�!�% "�%"�%"�%"�%"�%"�%"�%"�% "�%$"�%("�%,"�%0"�%4"�%8"�%<"�%@"�%D"�%H"�%L"�%P"�%T"�%X"�%\"�%`"�%d"�%h"�%l"�%p"�%t"�%x"�%|"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�%�"�% #�%#�%#�%#�%#�%#�%#�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍M�黽���T$�B�J�3��k����`��3���������������̡��������ËT$�B�J�3��5��������������������������������̍M��K����T$�B�J�3������� ��ö��������������̋T$�B�J�3��ӿ�����零����������������������̍M������T$�B�J�3�蛿������c���������������̍M�黼���T$�B�J�3��k�������3������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������|���h��������_^[���   ;�葟����]������������������������U����   SVW��@����0   ������j � ��2���_^[���   ;��<�����]������������������̋�U��Q3��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������	���_^[���   ;��Ύ����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �P���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            <%�B>A�K�,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            y)�%                                                                                                                                                                                                                                                                    }9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        z��O       o   $� $�	 IDM_NEU     SDK Test    IDS_EDITOR_PLUGINS      PLUGIN_CMD_1000472      M_EDITOR    C4DSDK - Edit Image Hook:       -plugincrash    -SDK executed:-)       -SDK    -SDK is here :-)       -help   --help              Baking in Progress...Please Wait                  �?    Controller Object_      Frame#           @�@    STEPS   tquicksteps     myicon.PNG          c:\program files\maxon\cinema 4d r12\plugins\quicksteps\source\quicksteps.cpp                   ���%B$V$"�@{6�="D+E�:�E~=47fK�A�'�-_C�5zF                    ܳ�L�?V$"�@Z%�="D+E�:�E�.47fK�A�'�-_CBzF                    ���:�?V$"�@Z%�="D+E�:�E�.47fK�A�'�-                %s(%d): %s      c:\program files\maxon\cinema 4d r12\resource\_api\ge_dynamicarray.h                i >= 0 && i < count     FALSE       c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp                 #   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp                %s      c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h                      �?             @�@          4&�k�          4&�kC        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basetime.cpp                      �Ngm��C           ����A        ����MbP?        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_memory.cpp               res �!E    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp                c:\program files\maxon\cinema 4d r12\resource\_api\c4d_string.cpp               no baselist      B   KB  MB           �@     GB c:\program files\maxon\cinema 4d r12\resource\_api\c4d_customdatatype.cpp               $��0�;I�DIJ�"�3gE^I        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp               ���1    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp                 شvE    t��;    ��qE    �	I    c:\program files\maxon\cinema 4d r12\resource\_api\ge_sort.cpp              �/      �?      �?3      3            �      0C       �       ��                              <�.        f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c            f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c                     fmod         to�C�C�CTC�C�C�C�C�C�C�C�C�C�C�C                                Unknown Runtime Check Error
       Stack memory around _alloca was corrupted
         A local variable was used before it was initialized
           Stack memory was corrupted
        A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                (�����l�8��                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                  Run-Time Check Failure #%d - %s         Unknown Module Name     Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s                   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                           Stack corrupted near unknown variable               Stack area around _alloca memory reserved by this function is corrupted
                %s%s%s%s    >   
   %s%s%p%s%ld%s%d%s           Stack area around _alloca memory reserved by this function is corrupted                 
Address: 0x    
Size:      
Allocation number within this function:            
Data: <    wsprintfA   u s e r 3 2 . d l l         %.2X    A variable is being used without being initialized.             Stack around _alloca corrupted          Local variable used before initialization           Stack memory corruption     Cast to smaller type causing loss of data           Stack pointer corruption        ��t�X�$���    f:\dd\vctools\crt_bld\self_x86\crt\prebuild\misc\i386\chkesp.c                  The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                       _ s e t d e f a u l t p r e c i s i o n                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c                         s i z e I n B y t e s   >   0           _ c f t o e _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c                         b u f   ! =   N U L L       e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                           _ c f t o e 2 _ l           s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o a _ l         _ c f t o f _ l         _ c f t o f 2 _ l       _ c f t o g _ l                   �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��                    tan cos sin modf    floor   ceil    atan    exp10   acos    asin    pow exp log10   log     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p                             p N o d e - > _ N e x t   ! =   N U L L                 s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                 f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c           FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    K E R N E L 3 2 . D L L         Client  Ignore  CRT Normal  Free    ����������    Error: memory allocation: bad memory block type.
           Invalid allocation size: %Iu bytes.
        Client hook allocation failure.
        Client hook allocation failure at file %hs line %d.
            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c                         _ C r t C h e c k M e m o r y ( )           _ p F i r s t B l o c k   = =   p O l d B l o c k               _ p L a s t B l o c k   = =   p O l d B l o c k             f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       Error: possible heap corruption at or near 0x%p                 p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Client hook re-allocation failure.
         Client hook re-allocation failure at file %hs line %d.
             _ e x p a n d _ d b g       p U s e r D a t a   ! =   N U L L           _ p F i r s t B l o c k   = =   p H e a d           _ p L a s t B l o c k   = =   p H e a d             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                                 HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()                _ m s i z e _ d b g         %hs located at 0x%p is %Iu bytes long.
             %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
                   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 DAMAGED     _heapchk fails with unknown return value!
          _heapchk fails with _HEAPBADPTR.
       _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADBEGIN.
         _ C r t S e t D b g F l a g             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t D o F o r A l l C l i e n t O b j e c t s               p f n   ! =   N U L L       Bad memory block found at 0x%p.
        Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              _ C r t M e m C h e c k p o i n t           s t a t e   ! =   N U L L           n e w S t a t e   ! =   N U L L         o l d S t a t e   ! =   N U L L         _ C r t M e m D i f f e r e n c e           Object dump complete.
      crt block at 0x%p, subtype %x, %Iu bytes long.
             normal block at 0x%p, %Iu bytes long.
          client block at 0x%p, subtype %x, %Iu bytes long.
              {%ld}   %hs(%d) :       #File Error#(%d) :      Dumping objects ->
      Data: <%s> %s
     ( * _ e r r n o ( ) )       _ p r i n t M e m B l o c k D a t a             Detected memory leaks!
     Total allocations: %Id bytes.
          Largest number used: %Id bytes.
        %Id bytes in %Id %hs Blocks.
       _ C r t M e m D u m p S t a t i s t i c s           o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g               Damage before 0x%p which was allocated by aligned routine
                  The block at 0x%p was not allocated by _aligned routines, use realloc()                 The block at 0x%p was not allocated by _aligned routines, use free()                _ a l i g n e d _ m s i z e _ d b g             m e m b l o c k   ! =   N U L L         CorExitProcess      m s c o r e e . d l l       _ w p g m p t r   ! =   N U L L         _ g e t _ w p g m p t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 d a t . c                         p V a l u e   ! =   N U L L         _ p g m p t r   ! =   N U L L           _ g e t _ p g m p t r       f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c             s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               _ s e t e n v p             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c            f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c            f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c          f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h e a p i n i t . c                       _ c r t h e a p           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                                      ��P�        ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                 _ v s n p r i n t f _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c                       ( f o r m a t   ! =   N U L L )         _nextafter      _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                �������             ��      �@      �                               ���5�h!����?      �?          r u n t i m e   e r r o r            
     T L O S S   e r r o r  
           S I N G   e r r o r  
         D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                            X   �	   �
   (   �   H   �
   �
   
   �	   0	   �   X          �!   Hx   $y   z   ��   ��   �                                        M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             
 
     w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                               . . .       w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           < p r o g r a m   n a m e   u n k n o w n >             w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                             R u n t i m e   E r r o r ! 
 
 P r o g r a m :                     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     _ N M S G _ W R I T E           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c                         s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         _ _ g e t l o c a l e i n f o               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t h e l p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\inithelp.c           M S P D B 1 0 0 . D L L     M S V C R 1 0 0 D . d l l               r   PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y                 S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S                       RegCloseKey     RegQueryValueExW    RegOpenKeyExW   A D V A P I 3 2 . D L L         D L L       M S P D B 1 0 0         ... Assertion Failed    Error   Warning     PH4    f:\dd\vctools\crt_bld\self_x86\crt\src\dbgrpt.c             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       p f n N e w H o o k   ! =   N U L L             _ C r t S e t R e p o r t H o o k 2                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c                           m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           Microsoft Visual C++ Debug Library          _CrtDbgReport: String too long or IO Error          s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                     Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)                    
Module:    
File:      
Line:      

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.                              m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                 <program name unknown>      s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         _ _ c r t M e s s a g e W i n d o w A           A s s e r t i o n   F a i l e d         E r r o r       W a r n i n g       ���    _ C r t S e t R e p o r t H o o k W 2           M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y                     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )                                     
 M o d u l e :         
 F i l e :         
 L i n e :         E x p r e s s i o n :               
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                     w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       _ _ c r t M e s s a g e W i n d o w W           _ c o n t r o l f p _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c                           ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c                       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )                                                                                         H H : m m : s s         d d d d ,   M M M M   d d ,   y y y y           M M / d d / y y         P M     A M     D e c e m b e r         N o v e m b e r         O c t o b e r       S e p t e m b e r       A u g u s t     J u l y     J u n e     A p r i l       M a r c h       F e b r u a r y         J a n u a r y       D e c       N o v       O c t       S e p       A u g       J u l       J u n       M a y       A p r       M a r       F e b       J a n       S a t u r d a y         F r i d a y     T h u r s d a y         W e d n e s d a y       T u e s d a y       M o n d a y     S u n d a y     S a t       F r i       T h u       W e d       T u e       M o n       S u n       HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun p f l t   ! =   N U L L             s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           _ f p t o s t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c                       _ g e t _ e r r n o             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d o s m a p . c                       _ g e t _ d o s e r r n o           s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                     _ f l t o u t 2             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c                         _ s e t _ o u t p u t _ f o r m a t             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t f o r m a t . c                               ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                   ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               B u f f e r   i s   t o o   s m a l l           ( ( ( _ S r c ) ) )   ! =   N U L L             s t r c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                     f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c           Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete      new    __unaligned     __restrict      __ptr64     __eabi  __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(    �5�5t5h5X5H5<545(555+� 5�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4|4x4t4p4l4h4d4`4\4X4T4P4D484,4 44�3�3�3�3t3P3,3 3�2�2�2`2@2,2(2 22�1�1�1�1�1t1D11�0�0�0l0@00�/�/+��/x/`/<//                                                                                CV:     ::  '   `   generic-type-   template-parameter-     ''  `anonymous namespace'       `non-type-template-parameter        `template-parameter     void    NULL    extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{        }'  }'  )   void    std::nullptr_t      volatile    ,<ellipsis>     ,...    <ellipsis>       throw(      volatile   const   signed      unsigned    UNKNOWN     __w64   wchar_t     <unknown>   __int128    __int64     __int32     __int16     __int8  bool    double  long    float   long    int short   char    enum    cointerface     coclass     class   struct      union   `unknown ecsu'      int     short   char    const   volatile    cli::pin_ptr<   cli::array<     )[  {flat}  s   {for    �;�;�;    �F� �=    �G0J�H    15�G�F    �6�)�(     ??     L8+�F    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h a n d l e r . c p p                         p n h   = =   0         _ e x p a n d _ b a s e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c                       p B l o c k   ! =   N U L L         ( s t r i n g   ! =   N U L L )         s p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c                         ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6             s i g n a l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c                       ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f:\dd\vctools\crt_bld\self_x86\crt\src\winsig.c             r a i s e       SystemFunction036           ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       r a n d _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r a n d _ s . c                       _ R a n d o m V a l u e   ! =   N U L L             ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c                         s t r   ! =   N U L L       ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c             ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 ( c h   ! =   _ T ( ' \ 0 ' ) )         (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       _ o u t p u t _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c                       ( s t r e a m   ! =   N U L L )         _ s e t _ e r r o r _ m o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c                         ( " I n v a l i d   e r r o r _ m o d e " ,   0 )               GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L             ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               w c s c a t _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                     w c s n c p y _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l                         w c s c p y _ s         s t r n c p y _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h                           ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                   _ w m a k e p a t h _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t m a k e p a t h _ s . i n l                         ( L " I n v a l i d   p a r a m e t e r " ,   0 )               _ w s p l i t p a t h _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t s p l i t p a t h _ s . i n l                           ( ( ( _ P a t h ) ) )   ! =   N U L L           f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t M o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c                         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   _ C r t S e t R e p o r t F i l e               _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       %s(%d) : %s         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed!       Assertion failed:           s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   , Line      <file unknown>      Second Chance Assertion Failed: File            _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t A           w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               _CrtDbgReport: String too long or Invalid characters in String                  s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       % s ( % d )   :   % s       w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                 w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d !           A s s e r t i o n   f a i l e d :                   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 
   ,   L i n e         < f i l e   u n k n o w n >             S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t W           GetUserObjectInformationA       MessageBoxA     s i z e I n B y t e s   > =   c o u n t             s r c   ! =   N U L L       m e m c p y _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c                       d s t   ! =   N U L L       _ s w p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s w p r i n t f . c                            _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                         _ s e t _ c o n t r o l f p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                             LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL  �^    �$�^L��K�^L��)�^L��3�^L�8�^L�6+                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         _ c o n f i g t h r e a d l o c a l e           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t l o c a l . c                       ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                       f:\dd\vctools\crt_bld\self_x86\crt\src\setlocal.c           s e t l o c a l e       L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     s t r n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ s e t l o c a l e _ n o l o c k           ;   =;  s t r c p y _ s ( p c h   +   s i z e o f ( i n t ) ,   c c h   -   s i z e o f ( i n t ) ,   l c t e m p )                         _ s e t l o c a l e _ s e t _ c a t             s t r c a t _ s ( p c h ,   c c h ,   " ; " )               _ s e t l o c a l e _ g e t _ a l l             s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   s t r n c p y _ s ( c a c h e i n ,   c a c h e i n S i z e ,   s o u r c e ,   c h a r a c t e r s I n S o u r c e   +   1 )                               C   s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   " C " )                 _ e x p a n d l o c a l e           s t r c a t _ s ( o u t s t r ,   s i z e I n B y t e s ,   (   * ( c h a r   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                           _ s t r c a t s             s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                               s t r n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   l o c a l e ,   l e n )                                             s t r n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                           _., s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & l o c a l e [ 1 ] ,   1 6 - 1 )                                             _ _ l c _ s t r t o l c         .   _   s t r c p y _ s ( l o c a l e ,   s i z e I n B y t e s ,   ( c h a r   * ) n a m e s - > s z L a n g u a g e )                         _ _ l c _ l c t o s t r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t t i m e . c                       p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                   f:\dd\vctools\crt_bld\self_x86\crt\src\inittime.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t n u m . c                         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initnum.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t m o n . c                         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initmon.c                                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                            _ _ s t r g t o l d 1 2 _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l                             _ L o c a l e   ! =   N U L L           1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 $ I 1 0 _ O U T P U T       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c                             _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r           _ v s n p r i n t f _ h e l p e r           ( " B u f f e r   t o o   s m a l l " ,   0 )               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   _ v s p r i n t f _ s _ l           f o r m a t   ! =   N U L L         _ v s n p r i n t f _ s _ l         ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   ( _ o s f i l e ( f h )   &   F O P E N )           _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c                       ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c                     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )               ( ( c n t   &   1 )   = =   0 )         _ w r i t e _ n o l o c k           ( b u f   ! =   N U L L )           f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c                         _ i s a t t y           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c          _ f i l e n o       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c                       p r i n t f         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p r i n t f . c                       _ w c t o m b _ s _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c                       s i z e I n B y t e s   < =   I N T _ M A X             _ m b s t o w c s _ l _ h e l p e r                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c                       s   ! =   N U L L       r e t s i z e   < =   s i z e I n W o r d s             b u f f e r S i z e   < =   I N T _ M A X           _ m b s t o w c s _ s _ l           ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                               s t r c a t _ s         l e n g t h   <   s i z e I n T C h a r s           2   < =   r a d i x   & &   r a d i x   < =   3 6               s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   s i z e I n T C h a r s   >   0         x t o a _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c                       x 6 4 t o a _ s         _ w c s t o m b s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c                       p w c s   ! =   N U L L         s i z e I n B y t e s   >   r e t s i z e           _ w c s t o m b s _ s _ l           ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               _ v s w p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c                       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s w p r i n t f _ s _ l         _ v s n w p r i n t f _ s _ l           x t o w _ s     x 6 4 t o w _ s         _ w o u t p u t _ l         _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             p l o c i - > c t y p e 1 _ r e f c o u n t   >   0                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t c t y p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\initctyp.c           united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american    D�ENU 0�ENU �ENU �ENA  �NLB ��ENC �ZHH �ZHI ��CHS ̐ZHH ��CHS ��ZHI ��CHT t�NLB `�ENU P�ENA <�ENL ,�ENC �ENB �ENI ��ENJ ��ENZ ďENS ��ENT ��ENG ��ENU t�ENU `�FRB L�FRC 4�FRL $�FRS �DEA ��DEC ��DEL ЎDES ��ENI ��ITS ��NOR ��NOR x�NON \�PTB D�ESS 0�ESB  �ESL �ESO �ESC ԍESD ��ESF ��ESE ��ESG |�ESH h�ESM T�ESN <�ESI (�ESA �ESZ �ESR �ESU ،ESY ��ESV ��SVF ��DES ��ENG ��ENU ��ENU                                                                                                         ��USA ��GBR x�CHN p�CZE d�GBR T�GBR H�NLD <�HKG ,�NZL (�NZL �CHN �CHN  �PRI ��SVK �ZAF ؋KOR ȋZAF ��KOR ��TTO ��GBR ��GBR |�USA ��USA                                     6-    Norwegian-Nynorsk           s t r c p y _ s ( l p O u t S t r - > s z L a n g u a g e ,   ( s i z e o f ( l p O u t S t r - > s z L a n g u a g e )   /   s i z e o f ( l p O u t S t r - > s z L a n g u a g e [ 0 ] ) ) ,   " N o r w e g i a n - N y n o r s k " )                                                   _ _ g e t _ q u a l i f i e d _ l o c a l e                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t q l o c . c                         OCP ACP #Cbad exception   ���3�G        i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                   s t r t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o l . c                       n p t r   ! =   N U L L         s t r t o x q       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o q . c                           ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 _ o u t p u t _ p _ l           ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f:\dd\vctools\crt_bld\self_x86\crt\src\osfinfo.c            _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c                           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                             f:\dd\vctools\crt_bld\self_x86\crt\src\_sftbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ s f t b u f . c                         f l a g   = =   0   | |   f l a g   = =   1             v p r i n t f _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v p r i n t f . c                         _ w o u t p u t _ s _ l         _ w o u t p u t _ p _ l         f p u t w c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t w c . c                       ( s t r   ! =   N U L L )           _ s t r i c m p _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r i c m p . c                         _ s t r i c m p         c o u n t   < =   I N T _ M A X         _ s t r n i c m p _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c m p . c                       _ s t r n i c m p       csm�               �                0�w5�G    Unknown exception       H��1�G    ���#�G     ��#�G    C O N O U T $       f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c                       _ f c l o s e _ n o l o c k         ( _ o s f i l e ( f i l e d e s )   &   F O P E N )             _ c o m m i t           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c                           ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         w c s t o x l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o l . c                       _ c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c                     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c                       s t r e a m   ! =   N U L L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 RSDSG,�0��K����x�L�   C:\Program Files\MAXON\CINEMA 4D R12\plugins\QuickSteps\obj\QuickSteps_Win32_Debug.pdb                                                                                                                                                                                                                                                                                                       �Ĳ               ز    ��X���     �       ����    @   Ĳ         �       ����    @   4�                   H�    �X���    <�       ����    @   |�                   ��    X���    X�        ����    @   ��                   Գ    ��                 �4�                <�|�                X���                ��<�               P�    \���    ��       ����    @   <�                    ����               ��    ��    ��        ����    @   ��                    ��               �    �4�    �       ����    @   �        4�        ����    @   X�                   l�    4�                4�X�                X���               ��    ��    X�        ����    @   ��                    x���               �    �    x�        ����    @   ��                    ��T�               h�    p�    ��        ����    @   T�                    ����               ��    ̶�    ��       ����    @   ��        ��        ����    @   �                   (�    �                ���                �`�               t�    ���    �       ����    @   `�                    8���               з    ܷ�    8�       ����    @   ��                    \��               ,�    <�ܷ�    \�       ����    @   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.�.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            .......................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ����    ����    ����    Wg    ����    ����    ����ej�j    ����    ����    ����    {k    ����    ����    �����u�u    ����    ����    ����FvLv    ����    ����    ����    ˭    ����    ����    ����    ��    ����    ����    ����    .�    ����    ����    ����    u�    ����    ����    ����    ��    ����    ����    ����    �����    9�        ����    ����    ����    (�����    ��        ����    ����    ����    <�    ����    ����    ����    ��    ����    ����    ����    M�    ����    ����    ����    1�    ����    ����    ����    v�    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    @�    ����    ����    ����    ;�    ����    ����    ����    ��    ����    ����    ����    .    ����    ����    ����=G=    ����    ����    ����    �X    ����    ����    ����    b    ����    ����    ����    A|    ����    ����    ����    �~    ������"�   X�                           ����    ����    ����    ��    ����    ����    ����    ��    ����    x���    ����    ��    ����    x���    ����    C�    ������"�   �                           ����    ����    �����~	�~	    ����    ����    �����	�	    ����    ����    ����m�	s�	    ����    ����    ����    ��	    ����    ����    ����    9�	    ����    ����    ����    �	    ���� �"�   ��                           ����    ����    ����    ��	        ��	        ����    |��    ����    7�	        ��	        ����    ����    ����    �	
    ����    ����    ����    �

����    
        ����    ����    ����    b
����    �
        ����    ����    ����    G
        L
        
            ����    ����    ����    �
    ����    ����    ����    �
    ����    ����    ����    ��
        �<    ��       ����        ��    ����       $        ��    ����       �D        ����    ����    ����    }M    MMZM        ����    ����    ����    �P    �OP        ����    ����    ����&U,U    ����    ����    �����V�V    ����    ����    �����W�W    ����    ����    ����{_�_    ����    ����    ����`,`    ����    ����    �����`�`    ����    ����    ����haua    @           �b����    ����                  P�"�   `�   p�                       ������"�   ��                           ������"�   ��                           ����    ����    ����    ��        s�        ����    ����    ����    3�    ����    ����    ����    ��    ����    ����    ����    "�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��        ��        ����    ����    ����    ��    ����    ����    ����    �Z    ����    ����    ����    �o    ����    ����    ����    5s    ����    ����    ����    ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        z��O    2�          (� ,� 0� �, A�   QuickSteps.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                       �    .?AVQuickSteps@@        �    .?AVTagData@@       �    .?AVNodeData@@      �    .?AVBaseData@@      8   Y  �  @     (   2   �   �   Q         v   �    .?AVResourceDataTypeClass@@         �   �   �  �  �    .?AVGeToolDynArray@@        -   �    .?AVGeToolDynArraySort@@        �    .?AVGeSortAndSearch@@       �    .?AVGeToolList2D@@      �    .?AVGeToolNode2D@@      �       u�  s�          �    .?AVtype_info@@         N�@���D                           �0�0�0�0�0�0�0�0�0�0        ?  ��������       ����   ��������    �����
                                                                             \�   X�   h�   `�   ,   $!      P�   H�   8�         �   �    �   0�   (�       �   �   �   �   �   �"   �#   �$   �%   �&   �                                                      �      ���������              �               �D        � 0                    0<                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                      ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ����C    ))))))) )�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(x(p(h(�(`(X(P(D(8(,( ((((�'�'	         �'�'�'�'�'�'�'�'t'`'H'0' ''�&�&�&�&�&�&�&�&�&�&�&x&d&L&<&,&�& &&&�%�%�%�%�%�%�%P%8%                                                                                                                                                                   L�            L�            L�            L�            L�                              ��        �o(t�uP�                                             � � �                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                         �&                                                                                                                                                                                                                                                                                                                                                               l1            �A�A    ����         ������������        �q    .   .   ��P�P�P�P�P�P�P�P�P���T�T�T�T�T�T�T���                    �o�q       ���5      @   �  �   ����                          �                    �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                  �    .?AVbad_exception@std@@         �    .?AVexception@std@@                      �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                            �    .?AVbad_cast@std@@      �    .?AVbad_typeid@std@@        �    .?AV__non_rtti_object@std@@         ����                                                                                                                                                                                                                                                                                                                                                                                    (          d) �!                     �# �# �# �# �# �# �# $ "$ .$ @$ P$ l$ x$ �$ �$ �$ �$ �$ �$ �$ % % &% 6% D% V% f% �% �% �% �% �% �% & & ,& F& V& l& �& �& �& �& �& �& 
' ' (' 4' F' V' d' n' z' �' �' �' �' �' �' �' �' ( .( D( Z( j( �( �( �( �( �( �( �( �( ) $) 4) B) P)                                                                                                             �# �# �# �# �# �# �# $ "$ .$ @$ P$ l$ x$ �$ �$ �$ �$ �$ �$ �$ % % &% 6% D% V% f% �% �% �% �% �% �% & & ,& F& V& l& �& �& �& �& �& �& 
' ' (' 4' F' V' d' n' z' �' �' �' �' �' �' �' �' ( .( D( Z( j( �( �( �( �( �( �( �( �( ) $) 4) B) P)                                                                                                             �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer WideCharToMultiByte  IsDebuggerPresent gMultiByteToWideChar �RaiseException  MlstrlenA  EGetProcAddress  ?LoadLibraryW  IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  GetLastError  �InterlockedDecrement  �GetCurrentThread  �HeapValidate  �IsBadReadPtr  ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter GetModuleFileNameW  %WriteFile GetLocaleInfoW  �HeapFree  �HeapAlloc JGetProcessHeap  �VirtualQuery  bFreeLibrary hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage � EnterCriticalSection  9LeaveCriticalSection   FatalAppExitA RtlUnwind �HeapReAlloc �HeapSize  �HeapQueryInformation  -SetConsoleCtrlHandler �InterlockedExchange �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -LCMapStringW  iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  GetLocaleInfoA  IsValidLocale EnumSystemLocalesA  �GetUserDefaultLCID  �SetStdHandle  � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 p (   p::�:;S;�;�;7<�<==�=>�>�?   � @   "0�01�122 2*23q3�3�3�34:4�46(646�6�6�78�9�:�:;   � 4   1Y5�5�5�5�6[7}7�7 8�8�8 99k9�9�;�;�;�<)>+? � H   0Y1�2�2�2�2 33-5�5?6�6?7�7@9h9t9�9:�:+;�;�;<g<�<�<�=�=`>0?   � P   �0�1�1�1�1j2�2�2�23�5}7�7�7�7�7�7�78H;W<a<f<s<�<�<�<=5???D?Q?t?�?�?�? � (   �3m4�4�5�67�7{8�8�9+;�;+<�<C>   � d   -020;0�0n1!2�2�23s3�3�3s4�4�4�4;5�5/6�6�6<7�7�788�8�8L9�9k:�:�:�:c;x;�;�<=�=�=�=�=�>;?   � X   k0�0�0�0�0�1;2�2Q3�4�4�4�4�4�5�6�6�6�6�67�7�7C8�8�8s9�9#:E:�:O;�;K<�<+=�=?>�>b? � P   {0�0_1�1_2�2_3�34<4H4�4/5�526�67�78o8�8n9�9[:�:O;�;R<�<4=�=>�>�>k?�?   @   K0�0+1�12�8�89�9�9�9�9_:�:�;�;�;q<�<�<f=k=y=>8>D>�>B?  L   L0�0,1�122�2o3�3O4�4_5�5O6�6(7�78�8E9�98:�:$;�;<t<�<_=�=m>�>F?�?   L   -0�01z1�1V2�3�3�364�4&5�56�6�6�78�8�8�9:�:w;�;T<�<;=�=>�>�>k?�? 0 P   K0�0+1�12{2�2[3�3;4�45�56�67�728�8<9�9:�:�:k;�;_<�<O=�=;>�>?�?�?   @ L   k0�0K1�172�23�3'4�45�5�5k6�6T7�7D8�8$9�9":�::;�;<�<�<h=�=r>�>_?�? P X   �01�12�23�34�4
5z5�5V6�6>7q7�7�7�7Z8�89�9�9f:�:m;�;?<�<6=�=>D>h>�>�>�>f?�? ` X   ?0�0�0f1�1M2�223�34�4�4�4�4Z5�5B6�67�7�7m8�8989D9�9:}:*;�;-<�<=}=�=]>�>:?�? p d   0�0111T1`1l1x1�1!2D2P2\2h2�2343@3L3X3�3c4S5?6�6K7�7K8�8/9�9:�:�:O;�;&<�<=�=>�>�?�?�?   � \   J0�001�1M2�2F3�3B4�4[5�5�6�6$7*7P7�7�7+808�8I9;:`:l:H;l;x;X<|<�<_=�=�=�=�>�> ?y?�?   � T   i0�0V1�1=2�23�3�3n4�4O5�5F6�6*7�78}8�8V9�96:�:;o;�;O<�<O=t=�=�=_>&?�?�?   � L   o0�0[1�1K2{23�3�3r4�4H5�5o6�6k7�7K8�8?9�9K:�:+;�;<�<+=�=>�>?�?   � D   0�01{1�1_2�2R3�3Q4�4Q5[6�6�6�8v:�:�:;<<<H<I=l=x=�=�>?? � 8   60\0h0+1�12�24,484F5l5x5�6�6�6�7�7�7�;�?�?�?   � D   �0 112@2L2�56o6�687�7D8o89�9^:�:K;�;?<�<;=�=?o?�?�?�?�? � L   R1�1K2�2+3�34�4�4o5�5�56676[8�8[9�9K:�:>;�;K<Y=|=�=�=�>�>�>�>m?�? � @   J0�01�1�2�3�3�3�3
44,4585`5e5�6�6 7%7B8R8v8�89�9�>        �6`7   H   �1�1k2�2O3�3K4�4D5�5+6�67{7�7[8�8R9�9K:�:;;�;w<�<r=�=o>�>r?�? 0 H   �01�1$2�2�2m3�3?4�45�5�5p6�6`7�7O8�8�9T:�:?;�;*<�<P=�=<>�>?? @ \   00a0F1�1�1p2�203a3�3%4�4�465�56E6�67Z78#8j8o8�89I9�9�9&:�:;v;�;V<�<R=�=R>�>�?   P H   �2�23m7w7�7�7�7�7�7�7�7�7�7�7�7�7�788949@9,:�>�>�>E?R?_?�?   ` x   �0�1$2�243�344�4Z5�5;6�6[78�89�96:>:�:�:�:�:;; ;b;h;u;�;�;�;�;<<<@<D<H<L<P<�<!=&=7=o=>>f>s>�>�>�>�>k?�? p ,   F0l0�0�0?1�1$202�23h3�3�34\4�5/8   �    o34@4L4 �    F7�7b8g8>?�?�? � h   �0�4555#5-575A5K5U5_5i5s5}5�5�5�5�5�5�5�5�5�5�5�5�5�5	616T6`67r;�;�;�;�;�;�;�;�;</>�>?�?�? � H   h0�0w12�23�34�4'5�5'6�6?7�7c8�8K9�9R:�:K;�;+<�<=�=*>�>?$?-? � (   �3�3�3�3�4�4�7(8�8?9�92:�>�>�>     L   �3�3�3�4�4/5�5�5�5�5x6}6�6?7d7p7|7�7h8�8o9�9_:�:R;�;g<�<_=�={>�>_?�?      80�0^1O5�9 :::$:O;o<�>   $   )2.2F2-9T9`9�9�:;8;D;�;(<h= 0    3)8�8J<�<�=�?�?�?   @ P   �1�1�1�1�1�1�1�1�1�1�1�122222$2+22292x2�2�2�2{34�45�56{6�6r7�7r8 P T   v7{7�7�7�:�:�;�;�;�;�;�;�;�;�;�;�;�;<<<<<<!<%<W<c<�<�<�<g=�=�=�=�=>? ` �   �0j1�1�1�1�1�1�1�1�12=2D2H2L2P2T2X2\2`2�2�2�2�2�2"3-3H3O3T3X3\3}3�3�3�3�3�3�3�3�3�3�3F4L4P4T4X4�5(6-6?6�6�6�6�6�677!7.7_7�7�7�7�7�7999D9g9|9�9:@:U:(;-;?;�;�;�;�;S<�<�<�<�<�<�<�=�=�=�=�=>�>a?k?�?   p �   g1n1�1�1�1�1�1�1 2'2B2�2�2"3F3�3�3�34A4i4(5-5?5~5�5�5�5@6�6�67<7p7u7�7�788'8.838N8T8]8f8k8v8�8�8�8�8�8�8�9�9�9:B:|:�:�:@;c;j;�;�;�;�;�;�;�;�;<<<V<f<z<<�<Y>j>�>�>   � d   �1$202]2b2g2�2�2�2�2�2.4:4g4l4q4�4�4�4�4�4(545a5f5k5G6L6Q6V6K729>9k9p9u9�9�9�9�9�9&:2:_:d:i: � t   �23 3M3R3W3|3�3�3�3�355<5A5F5x5�5�5�5�5�7H8T8�8�8�8�8�8�8�8�8t<{<�<�<�<�<�<�<�=�=�=�=>>7>E>�>�>)?u?�?�? � �   0d0�0�091T1�1�1=2�2�2�2�2A3L3�3�3�34U4`4�4�45Y5�5�5J6�6�6�6 77777777 7$7(7,70747�7�7�7�7�7�7�7�7 8888�:�:�:;;>;�;�<�<�<�<�<2=<=�=�=8>=>O>u>z>7?<?A?   � �   H0M0_0�0�0�0�0�1�1�1�1�1l2�2�2 344/497W7{7�7�7�7�7�7�7�7�78&8I8O8i8s8x8}8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89
9999%9,9A9H9M9S9Z9_9e9l9q9v9}9�9�9�9�9�9�9�9�9�9�9 :�:�:�:�:�:�:�:�:;8;=;O;c;i;v;�;�;<�<�<�<�<�< ==J=�=�=�=�>�>?d?m? �   W0e0l0v0}0�0�0�0�0�0�0�0�01#1�2�2�2�2�233 363B3K3P3Y3e3n3�3�3�3�3�34k4p4�4�45*535;5D5L5R5X5`5f5l5t5�5�5�5�5�56899/9/:8:A:Q:]:s::�:�:�:�:�:�:�:;;E;f;�;�;�;<%<b<n<�<�<==�=�=�=�=�=�=�=�=�=�=�=�=>>>>>A>]>�>�> ?
??2?P?Z?f?�?�?�?�?�?�?   � �   h2m22�2�2�2�2�2�3�3�3x4�4�4�4�4�4�4�4�4
565Q5]5b5�5�5�5�56$6t6z6�6�6�6.747l7r7�7�7�78(8A8J8O8u88�8�8�8�8�8�8979�:�:�:�:;.;3;8;N;W;`;p;|;�;�;�;�;�;)<5<=#=H=M=_=�=�=g>s>�>�>�>?#?�?�?�?�?�?�?�?�?�?   � �   00E0�0�0�0101V1�1�12=2a2�2�283<3@3D3h4m44�4�4�45	55545K5a5g5t5666E6Q6~6�6�6�6�6�7�7�7�78�8::6:H:M:_:�:�:�:�:�:�:+;�;�;<&<==<=A=F=l=x=�=�=�=�=�=>>>�>�?�?�?   � �   0 0I0�0�0�0171�1�1�1�12]2�2�2�3�4�4�4�45	6,6<6A6�6�6�6�6�6-7I7m7�7n9z9�9�9�9�9�9(:-:2:�:9<V<�<�<�<�<===U=a=�=�=�=l>     �   �0�0 11�1�1�1�1N2Z2�2�2�2h3p3�3�3�3�3�3�3�3�3�3�45,555k5z5�5�5�5�5�5�5�5�5�5�5�5�56666�6�6�6�6�6�6�6�67
7p7�7�7�7�7�7�7�7�7�78D8�8�899W9�:�:;	;;%;7;C;p;u;z;�;�;<4<9<><U<g<s<�<�<�<�<=(=P=V=j=8>K>g>|>�>�>�>g?�?�?�?    �   :0[0�011V2c2{2�2�2�2
33l3�3�3�3�3
44.43484l4{4�4!5/5:5B5G5U5]5j5v5�566y6�:G;W;x;�;�;<<.<D<K<^<�<�<�<�<�<�<�<�<==]=>&>>>_>�>�?   �   000'0<0H0T0d0�0�0�1�1�1�3�3,42484>4D4J4Q4X4_4f4m4t4{4�4�4�4�4�4�4�4�4�4�4�4�4�4�4555&5�5�5�5�5�596B6l6q6v6�7s89m9O:�:#?�? 0 H   �0�0�0�0V3a3�3�3�3�3�3�3�4�7�7<'<<<�<�<�<�<�<�<L=�=�=8>�>D?�?�? @ �   �0�0�0�0�0�0y2�2�3�3�4�4505t5�5�56�6�6R7n7y7�7�7�7�7�7�7�7888m8r8w8~8�8�8�8�8�8�8�8�89"9'9:�:�:(;S;X;];�;<]<�<�=�=>`>i>v>�>�>�>�>�>�?�? P �   <0C0<1G1`1u1{1�1�1l2w2}2�2�2�2�2�2�233R3�3�3�3�3�3�3�34�4�45�5�5�5�56.63686_6h6�6�6�6�6Q7j7s7�7�7888Z8c8l8�8 :^:n:s:x:}:�:�:�:�:f;r;�;�;�;�;�;�;<<)<9<E<q<�<�<�<�<==D=I=N=�=�=�=�=�=??/?k?t?�?�?�?�?�?   ` �   00030�0�0�041l1u1�1�1�1�1�12�3�3�3�3�3�3H4M4R4Y4�4�45 5,5@5L5g5w5�5�5�5�5�5666*6�6�6�6�6�6�6�6 77,7-969`9e9j9�9:$:�:�:�:�;�;�;~<�<�<�<�<�<>�>�?   p \   �0�1�2g3W4G5767;x;};�;�;�;�;<<"</<�<�<�<3=�=�=�=�=>>>I>x>�>�>�>�>�>�>�>�>?   � h   00C0S0]0�0�0�0Y1�12T2�23%3l4�5�5�5�5�5�5�5�6�6,7E7�;�;�;<4<P<l<�<�<�<=v=�=�=�=�=>5>i>�>�> � p   W0�0?1K1�2(3-3?3b3�3)4�5	7�8�8�8�8�8�89/94999t9}9�9�9�9�9�9:::'<3<�<='=,=1=�=�=>>>u>�>�>(?-?2?   � �   Y1s1|1�1�1�1�1�112:2d2i2n2�2�2�2�2)3.333�3�3�344D4I4N4�4�49,969N9U9c9�9�9�9�9:-:::G:T:�:�:�:�:�:;M;_;�;;<b<i<�<�<�<�<�<�<;=k=�>�>�>�>,?�?�?�?�?�?�?�?   �   0000%0}0�0�0�0�0�0�0�01"11�1�1�1�1�1�1�1�1�12�2,393b3l3�3�3�3�3�3�3�3�3�34d4u4�4�4�4�4#5�5�5�5�5�51667D7h7q7�7�7�7�78!8F8O8X8c8l8q8�8�8�8�8�8�8�8�8�8�849S9`9�9�9�9�9�9:":5::;I;R;x;;�;�;<+<3<9<]<o<�<�<�<�<==%=K=R=X=a=y=�=�=�=�=�=�=)>4>K>V>�>�>�>?4?B?Q?Z?�?   �   �0�0�0�011#1H1P1i1�1�1�1�1222)242C2i2v2~2�23@3D3H3L3P3T3X3�3�3�3�3�3�3�3�3�3�3�3�3�3P4T4X4\4`4d4h4�6�6�67	77.777Y7e7s7|7�7�7�7�7�788I8\8g8�8�8�8�8�8'9.949C9Q9Y9�9�9�9�9�9$:5:P:c:p:y:;_;�;�;�;�;�;�<===�=�=�=�=�=�=�=>> >K>^>g>�>�>�>�>?5?=?H?P?X?   � �   �0111,151N1\1o1|1�1�1�1�1�1�1,2:2[2d2j2r2{2�2�2�2�2�2�253�3�3�3�3�3�3Y4s4�4�4�4�4�4�4	55'5/545G5T5c5l5�5�5�5�56*6l6z6�6�6|7�7�7�7�7�7�7�7�7�7$8U9�9�9�9�9�:7;@;p;t;x;|;�;�;�;�;�;�;�;�;�;�; � $   �0�0�45|6!7G7T7{9�:a;<D=V> � x   	0�0w1"2�2�2�8�8�8�8�8�8�89O:�:;;;3;:;�;�;�;�;�;�;�;�; <<<!<'<5<B<K<T<�<�<�<�<�<�<�<�<=)=�>�>�>�>�>�>�>?  	 �   ]1k1t1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1@2D2H2L2P2�2�2�2�2�2�2�2�2�2|5�5�5�5�5�5�6�6�6�6�6�6�6*7�7�7�7�7 8'8�8�8�8 99999�9�9�9�92:;:L:g:~:�:�:Q;k;r;�;�;�;�;�;<G<P<U<o<v<|<�<�<�<�<�<�<=J=S=Z=�=�=�=�=�= >>>>>X>\>`>d>h>l>p>t>x>�?�?�?�? 	 L  00'0,0]0�0�0�0�0�0�0�1�1�1�1�122)2G2U2h223&343=3m3�3�3
444U4\4a4s4�4�4�4�4�4�4�455&575I5[5m55�5�5�5�5�5686A6R6a6p6x6�6�6�67B7I7R7�7 858L8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 999h9l9p9t9�9�9Z;e;m;�;�;�;�;�;�;�;�;�;�;<t<x<|<�<�<�<�<�<�=�=�=�=�=�=>#>/>8>W>^>g>�>�>�>�>�>�>�>�>�>�><?c?p?~?�?�?�?�?�?�?�?    	 x   i0�0�0�0�01M2�4�4�4�4Q6Y6_6�6�6�6�6�6�67777'7_7n77�7�7�7�788#899^9g9�:�:�:B;K;s;�;�;\<z<�<�<==!=�=�= 0	 �   �1�1�1�1�12-2:2B22�2L3�3�3�4[6�6�6�7�7�7�7v8�8�8�89F9S9[9m9z9�9�9�9�9�:;2;@;I;�;F<f<�<�<�<�<=&=F=f=�=�=�=�=>">F>n>�>   @	    �29)9�: P	    �1D45�5+7�;>r>�?   `	 |   �0�0�1�1h3�475e5�5�5�5�5�5�5�5�56.656�6<9�9::N:U:d:�:�:�;Y<�<�<�<�<�<�<==7=>=�=�=�=�=>	>E>L>^>e>�>?"?�?�?�?   p	 �   	060�0�0/181b1g1l1�1�1�1�1�1�5�5�5�58#8�8�8�8�8�8�8�8�89?9]9d9h9l9p9t9x9|9�9�9�9�9�9�9B:M:h:o:t:x:|:�:�:�: ;;;;;;;;f;l;p;t;x;�=�=�=�=&?,?1?H?M?_?   �	 �   00/0F0M0�0�0�0�0111�1�1�1�1�1�1�1�1 2222&292>2F2M2`2e2m2t2�2�2�2�2�23$3�3�3�3�3�3*4/444\4`4d4h4l4�4�4�5�5�5�5�5�56�6�6�6777:7W7t7�7�7&8+808J8�8�8�8�9�9�9�9�9�9�:�:;;i;�;�;�;�;�;�;�;<<F<O<y<~<�<�<�<�<�<�<== =.=C=W=]=l= �	 `   82G2?3H3�4�4F5R5�67)7Y7^7c7�7�7:8L8�8�8�8�8�89&9V9[9`9:9:h:�:�:;;;�;�;�<�<> >�>�? �	 h   (0�0�0111�1s2z2�2�2�2�2d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9   �	 �   �01�1@2D2H2L2P2T2X2\2�23383A3k3p3u3�3�34$4*4?4I4c4h4m4w4~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4555o5z5�5�5�5�5�5�5�6�6�6�6�6C7K7�7�7�7�7�7<8D8q8�8�8�8�8�8Q9X9�9�9�9�9�9�9+:3:�;�;�;�;�;8<@<�<�<�<�<= =%=�=�=M>U>�>�>�>�>�>�>(?0?   �	 �   �0�0$1)1.1s1{1�1�1�1�1�1}2�2�2�2�2333W3_3�4�4�4�4�4&5.5�5�5�5�56	66}6�6+737^7�7�7�7�7�788�9Q:y:�:r;~;�;�;<<<F>N>�>�>�>??:???D?   �	 �   �1�1�2�2�3�344z4�4�4�4C5K5�5�5�5�5�5
66C6H6M6A8J8x8}8�8�8�8�8�899+9;9�9�9:::7:C:T:^:n:x:�:�:�:;;;6;�;<<<#<K<Q<l<y<~<�<�<�<�<=="=X=]=b=g=�=�=�=�=�=�=�=�=*>;>@>E>J>s>x>}>�>�>???S?X?]?b?�?�?�? �	 �   0
0070<0A0F0i0r0�01�1�122D2K2U2g2q2�2�2�233H5M5f53696M6R6W66�6�6�6�6�6�6�6�6B7G7L7�7�7�7�7�7�7�7�7�788 8T8e8j8o8t8�8�8�8�8	9=9B9G9}9�9�9�9�9�9�9�9 ::L:Q:V:[:~:�:�:0;�;�;<0<A<H<�<�<�<�<�<�<8=?=z=�=�=�=�=�=�=�=>>D> �	 �   �0�01
11)1C1H1M1W1^1c1h1r1y1~1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1O2Z2a2{2�2�2�2�2�3�3�3�3�3"4+4U4Z4_4�4�4�4�4�4�5�566"6I6U6�6�6�6;^;$<=/=8=�=�=�=�=  
 P   �7�7>8q8�8�8�8�8�8�8�8 99X9]9o9�9�9�9�9�9::/:o:}:�:�;!<i<�<�>�>�>�>�? 
 d   00/0y0�0�0�0�0�0�1�1�1�13"3(33393E3l34�4�4�4*5/545\8%9�9�9�9q;�;X<�<�<�<�>\?h?�?�?�?�?    
 h   0"0Y0o0�0�041J1|23333]4i4n4s4�4�4�4	666�6�6�67[7`7e7�7�7�7888�899;9j9�:%;M;�;+<U<�< 0
 (   �2�4�4�5�5�5�9P:o:�:Q;^;v;�;�;   P
 @   �3�34U5`5l5w5�5�5�5�5�568%8D8c8�89/9y9�<l=�=�=�=�=   `
 H   H0g0�0�0�0�01!1@1_1~1�1�1^2l2{2�2�2�23I3f;�;�<==J=O=T=�=?? p
 D   r0y0g1n14686<6@6D6H6L6P6T6X6\6`6d6h6l6p6�6�6�6�6�6 7�9:':	; �
 X   	1�1�2�2�2�20353:3?3�3�3�3�3�3�3�3�3�;<<�<�<�<_=h=�=�=�=�=�=�=�= >�?�?�?�?�?   �
 �   p0�0�01_1h1�1�1�1�1�1222�3�3b4n4�4�4�4�4�45 5%5N5�5�5�5�566"6`6g6�7�7�7�7�728>8k8p8u8�8�8�8k9�9�92:>:k:p:u:�:�:;<�<�<�<�<R=u=~=�=�=�=�=�=><>A>F>�>�>�>�? �
 �   060E0x0�0�0�01Q1t1}1�1�1�1�1�1282=2B2{2�2�2�3�3�32474<4b4�4�4�4�4�45F5�5�5�5606G6S6y6�6+7J7�78#8H8�8�8�89O9t9�:�:�:�;�;<2=G=�=�=�=>>7>�>   �
 �   �1�1�1�1�1�2�231363;3]3�3�3�3�3�3�3�3�34
44"40464f4o4�4�4�4�4]5n5�5�5�5�576X6a6}6�6�6)727\7a7f7�7�7�7�7�788"8):4:F:]:�:�:�:;/;4;9;�;�;<<<�<�<==5=:=?=�?�? �
 �   0!0&0�012�244�4�4�4�4�4(505�5�5�5�5�5]6d6�6 7=7I7v7{7�7!9*9T9Y9^9�9�9�9�9::#:�:�:�:�:�:$;);.;�;�;�;�;<2<7<<<|<�<K>T>~>�>�>�>�>�>�>�>#?+?n?w?�?�?�?�?�?   �
 t   0"0'0�0�0*1/141q3}3�3�3�3�3�3444U4]4�4�4�4�4�4"5.5[5`5e5[6g6�6�6�6)8f8o8�8�8�8�9Y:�:�:�<d?p?�?�?�?�?�?   �
 �   V0b0�0�0�0�01�1�1�1�1�1223�3�3�3�3�3484=4B4K6�677K7P7U7�7�7�7�7�7�788?8�8�8�8�8�899I:U:�:�:�:�:�:; ;%;g;�;�;!<�<�<�<�<'=,=1=q=y=?m?   �
 �   ;0D0n0s0x0�0�0�0�0�011b1k1�1�1�1�1�1222�2�2'3,313�5�5�5�5�5�5�5"6'6,6g6o6�6�6�6�6�667B7o7t7y7x8�8�8�8�8\:�:�:	;;;U;a;�;�;�;A<v<�<1=8=G>N>�?�?   l   f0/1�1b2n2�2�2�2�34464=4k4r4�9�9�9 :::::::: :$:(:@:D:H:L:P:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:    \   1+1X1]1b1�1�1�1�1�1�3�3(4-424�4505b5�56676R6m6�6949�:�:�:�:�:�:�<�<^=l=�=�=>,>   `   1�2�2�2�2�25:: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:p>�>�?�?   0 @   $0)0.030d0�0�2�23^3�3Q5�8�8�8N9;;\;�;�<�<=3=<=d=�=R> @ $   &0D0�3�3*8N8�8X<]<o<(?-???   P (   �2�2�2�5�56H7M7_78?=?O?�?�?�?   ` \   x0}0�011/1�2�23�3Y577h7w7�7�7�7�7�7Q8Z8�8�8�8�=�=G>]>�>�>�>?0?5?:?�?�?�?�?�?   p L   G5]5�8�9�9:::�:�:�:;J;V;�;�;�;�;�;<<<b=�=�>�>�>�>�>�?�?�?�?�? � �   40�0�0111�1�1�2	393>3C344@4p4u4z4�5�56"6'67$7T7Y7^7"8)8�9�97:C:s:x:}:G;S;�;�;�;�<�<�<�<�<�=�=�=�=�=�>�>???�?�?   � �   000�0�1�1222�2�2333�3	4�4�4555�5�566!6�6�6�6�67�7�7*8/848�8�8-92979�9�:�:�:�:�:;";�;�;�;�;%<,<�=�=�=�=�=�>�>�>�>�>�?�?   � t   000�0�0$1)1.12'2W2\2a2+373g3l3q3D4P4�4�4�4T5`5�5�5�5{6�6�6�6�6�7�7�7�7�7�8�8�8�8�8�9�9�9�9�9J?V?�?�?�?   � h   >0z1�1�1�1�1 2$2(2,2024282<2@2D2H2L2P2T2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2$3(3,3034383<3@3 � h   4�4�4�4�4�4V5h5�5�566>6C6H6�6�6�6�6�6t7�7�782878<8�8�894999>9�9�9�:;8<?<=�=G>�>�>*?/?4?   � p   0�0�0�0�0�0�0�6�6�6�6�6074787<7@7D7H7L7P7T7X7\7`7d7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7H?M?_?�?�?�? � �   E0�0�0�0�0%1+141I1�1�2�2�233"383�3�3�34(444@4V4�45&5^5c5h5�5�5�5�5�5�56�6�6�677�7�7�7�78K8i8H9M9_9�9�9::�:�:�:�:�:x;�;�;�;M<V<!=�=�>�>�>??.?D?m?z?�?�?   � �   80=0O0x2}2�2�2�2�2333O3y3�3�3�4�455-575V5�5C6O6�6�6�60797c7h7m7R8�8�8�89@9l9�9�9::#:e:q:�:�:�:Q;�;�;�;<<<d<�<�<>>A?H?   t   %0�0q1!2-2]2b2g2C3�3�3�3�3*414�9�9:	::\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;  \   �4�5�5�5�5�56)6Y6^6c6�7�799>9C9H9�9�9&:+:0:~:T;[;m<y<�<�<�<�=�=�=�=�=S?_?�?�?�?     �   �0�0�0�0�0�1�133�3�3�3�3�3�4�4�4�4�4A6M6}6�6�6S7_7�7�7�78@9L9|9�9�9R:^:�:�:�:;�;x<�<�<�<�<�=�=�=�=�=k>w>�>�>�>�?�?�?�?�? 0 �   �0�0�0�0�0�1K2W2�2�2�2�2�2]3d3�3�3�3�3[5g5�5�5�5m6y6�6�6�6�7�7�7�7�7�8�8�8�8�8�9�9:::�:�:%;*;/;<<><C<H<= =P=U=Z=;>G>w>|>�>M?Y?�?�?�?   @ �   c0o0�0�0�0u1�1�1�1�177B7G7L7�799N9S9X9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:::::H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�: P 8   (:-:?:e:n:�:�:�:i;�;�;4<@<==W?`?�?�?�?�?�?�?   ` �   00�1�12+20252^2g2�2�2�2Q3Z3�3�3�3�3�3�3�3474@4j4o4t4�56$6Q6V6[6�6�6�6�6�6�6�6)7.737�8�8�8n9�9�9�:�:�;j<�<�<:=^=�=
>.>e>k>p>�>�>�>�>�>�>�>�>?/?4?9? p �   "0+0U0Z0_0H1M1_1�1�1�1�1�1�1242=2g2l2q2�2�2�2
3394B4l4q4v4�4�4�4�4�4?9H9�:�:L;X;H=M=_=�=�=�=>>>2>J>S>�>�>�>�>?
?   � �    00M0`0�0�0�0|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 666666$6*60666<6B6H6N6T6Z6`6f6l6r6x6~6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777 7&7,72787>7D7J7P7V7\7�:�:�: ;:;b;�;�; �    <<q<   �    �<   � �   1114 4$4(4,4<7@7H8H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ??? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?   � p   22H3L3P3T3X3\3`3d3h3l3�3�30444<4@4H4L4T4X4�455�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�54989<9@9D9H9�=�=�=�=�= �    �7�7�7�7�7     8   �1�1�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>     \6`6d6�<�<�< 0 �   �5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777770;4;8;@;D;H;P;T;X;`;d;h;p;t;x;�;�;�;   P ,   �>�>�>�>�> ???????? ?$?(?,?   � �   P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4�6�6�6�6 �     �8�8�8�8�8�8�8�8�8�8�8 9 � @  �2�2�2�2�2�2�2�233(3@3H3L3P3X3p3�3�3�3�3�3�3�3�3�3 44440444H4P4T4\4t4�4�4�4�4�4�4�4�4�4555(545L5d5l5�5�5�5�5�5�5�5�5�5�566606H6L6`6h6p6�6�6�6�6�6�6�6�6�67 7(7<7@7T7X7l7t7x7�7�7�7�7�7�7�7�7�788$8,80848<8T8�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>   � �   �0�0�0�0�0�01101P1p1�1�1�1�1 2202P2p2�2�2�2�2303P3p3�3�3�3�3�3404P4\4h4�4�4�4 555L5P5l5p5�5�5�5�5�5�56@6L6p6|6�6�6�6�6�6 7,787`7�7�7�7�7�7�7�7�7�78(80848X8`8d8�8�8�8�8�8�8�8�899$9(9D9H9\9�9�9�9�9�9�9�9(:4:X:x:�:�:�:�:;(;H;h;�;�; � 8   0 0<0X0�0�0141X1x1�1�1�1 22222222�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�344H8P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;X<h<x<�<�<�<�<�<�<�<=== � H   P0`0d0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�011h1p1�4�4888\8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            