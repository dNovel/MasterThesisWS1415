MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       $�E�`�+�`�+�`�+��ӳ�a�+�{ ��w�+�{ ���+�i布c�+�`�*�1�+�{ ��&�+�{ ��a�+�{ ��a�+�Rich`�+�                        PE  L �u=P        � !
  �  �     [�                             �         @                   �8 `   � (                            � x:  `<                                            ؑ �                          .textbss=�                        �  �.text   ��  �  �                   `.rdata  P
  0    �             @  @.data   �B   @     �             @  �.idata  	   �     �             @  �.reloc  dD   �  F   �             @  B                                                                                                                                                                                                                                                                                                        ������� �!% �\� � �NG ��� �� �cr �nd �9~ ��e �� �� ��9 �pT �3 �f� ��# �<� �2 �r� ��I �(� �s� ��G  �x � ��) ���  饟 ��X � �&p �A�  �L �'� ��m �� �h �sJ ��5 �  �bG �/ �ZI �H � 髣 �VK �� ��h ��� �� �H  �rF �1 ��V �Y �D� �_9 �r �+F �P �+ �V� �1� �\ ��� ���  �-�  �  �3 �n ��� �� �oA ��  鵷 ��P 髧 ��= �q� �|, �ǐ �B� �}� ��  �7 �> ���  �� �= �  ��x ��  ��' ��@ �� �L^ �- �B� �0 ��� ��1 �Na �! �4+ �? �ڳ  �� 鰔 鋄 ��� �D �,u �/ �R# �� ��] �3 �  ��� 餀 �O�  �� 饔 � � ��  �V% � �~ �� ��z  �� �(� �C� �r  �Y; �tD �_� �z� ��� �� �^ ��1 �a 鬼 � �2 �m� �(R ��  �N� �9% �t�  ��C �d 饁  �P �ˁ �, �� �l� �- �b~  �M�  �H' �3�  �J 鹝 �d� ��� �� �J ��� �+� ��  �a�  �LB �w�  �r�  �]% �h� �cQ ��� �v  �4l ��  �� �� � � �+ �Fx �b �( �, �"� ��) �x�  �s� ���  �I� �4� �� �] �� �PC �K� �� �1J ��
 �� � �=� �� �S �~ �9 �_ �� �� ��b �r  �� ��� �* �H 鷁 �r' ��H  �+ �� ��� �[ ��E  �� �:� 饓 �[ �{� �v[ ���  �LC ��c �' �B �D ��� �G  �T �� 韃  �� �S � ��  �� ��� ��> ��[ ���  �� ��|  �� �� �YG �d�  ��A �zV ��� � I �+� �� �� �, �'� ��� �� �8) �S� �. �I� �o �OG �8 �u� �0( �+ �& �cA � �� �$A �m� �H2 �C ��B �	( �� �� �A �� � & �? ��j  �!C �\ �^ ��s �MT � 郮 ��� �Y�  ��� �] 銔 鵍 � �{G �6� �q� �� �G� � �m� �X� �� �� � �A ��F ��y �U� � �[% 鶨  �!
 �l 釞  ��  �]� �x�  �S �� �9 �$$ �?� �*� �� �� ��  ��P �& ��N �w6 �E �Ms �x�  �S� �^O ��� �:A �_H ��� �� �@I ��  �&� �( �G ��� �; �}� �� �c �  �I� 餹 �3 ���  鵁  �% � 鶏 ��� �^ �'� �� �}� �H� �L �N� �9�  �� �	 隩 �� �@" � ��? ��G �,R 駣 ��? �M' �H( �< �~4 �l �DF �- ��z �e@ �0' �� �� � ��  �'�  ��' �=� 鈎 �s�  ��( �9_ �$�  ��% �ʱ �U" �\? �� ��D ��U �,� � �i ��? � �� �~! �YD 锫 �� �
�  �5E ��� �k[ �� ��  � � �� ��< �X�  �s� � �? �� ��m �j ��Z �� �k� �6�  �� ��> �G� �Rm 鍥 ��� �CN ��  �ɸ �= ��m ���  �e[ �0  ��  �v� �� ��k  �> �� �M �(� �� ��Y 鹁  �d� �J �J �%^ �P�  ��� ��	 � ��  ��x  ��� �� � �� �.S �� 餯 ��� �� 镫 � �� �,= �ѹ �\ �G �? � 鸥 ���  �� �` �` ��� ��> �u� � � �B  �< �a �� �W� � �� ��= �c{ � �Y�  � > ��� 麍  ��� � �  �[ 醕  �Qp  �n  ��" � �� �} �s �>� �0 鴍 ��  �.? 饒 �`� 髷  �$ ��  �\� �w� �R �F �B �c�  �n� �� �4> � �
� �� �0� �� �' �y �\\ ���  �� �� ���  �S# �n� �y� �" �� �z�  ��  �� ��1 �6 �!� �,� � �2M �� �x �� �3 �	& �T� �+ �l; � ��� �k� �&� ��N ��  �'t  ��l  �}p �xw  �: �.� ���  �; �/ ��� ��� ��k  �k�  �x �� ��� �7A � � ��A �Cn ��� ��Y �TH �?�  �j�  �5 �Ъ �K� �VW �Q' 錉 ��A �b �� �) �# �H �yB ��� �o� �*� �E� �+ ��K �&d �� �@: �o �r� 魺 �� ��: �� �y� �D �/� �J) �5) �m  �k� � �! �� �� �) ��� ��' �S�  �>�  �	j  餾 �/� �:� ��x �  �' �2 �� 鼰  �ף  ��g ��� �T ��  �N� �y� �4v  � �J� 酠 ���  �K� ��� �!\ �� ��H ��  �j �X� ��  ��  �y< � �> �z: �5- � K �+� �6� ��S �� �� 邡 �M� �� �#w �/ �9  ��;  ��  �: ��
 鰱 �� ��� �9 �8 駂 �b2 �-�  ���  �l �n� �Y{ 餃  �; � �e�  �8 �� � � �� �G� ��? �� �� �� �~� ��  鄪 � �* 饪 �а �� �F�  �q� �O 釸 �29 �? �8 �� �^n �� �t�  � �j�  �5 � �;� �6; �q� �"9 �� �@ ��� �} �� �N�  �i7 �t� �� �jt �; ��W ��  �< �E7 �<m 駤 �a �}� �h�  �c_  �� �y�  �; �8 銦 �� �Y ��� � �� �L �H �¢ ���  ��{ 链 �N^ � �$A �� �V �� �Ћ ��6 ��� ��� �4 �'� �� ��� ��~ �e  �n� �I� �~ ��5 ��� �" ��A �{� � �F �� �G� �� � 鈬 �s� �>+ �iI �� � ��) �e� � � �x ��  �a�  �L�  駭  � �� �ؤ �� �� �i" ��� ��f � �E; ��:  ��/ �j ��� ��5 �( �R> �� �x� �s�  ��( � �,7 �O� �:�  �%; �`7 黒 �& �� ��i  鷻 �RQ ���  �x� ��  �>o �� ��= �O� ��  �u� 逖 ��$ �V�  �1� �,D �w� � �� � �c� �> �9� ��T �G �J� ���  �`�  �KF �&�  �ч  �L�  �G` �"� �� �� �� ��  �� �� �_h � �E� � L �+^ �& �Q �lm � �"� �Mp �� �c* �n� �� �* �H �JY �5 �п �� ��8 � �< �� �� �ͤ ��� �} ��� �9� �T* �_a ��& ��m  �`6 �k �6�  鱿 �} ��W �r�  �| �ȅ �� �.1 �9�  �� �/# �z ��r �`> �4 �f� �q�  �l�  �gP �b �M �4 �c ��� ��� �$� 鿜 �J5  �A 頞 ���  �y �a �,� �ט ��� ��6 �hR ���  �^�  �� �$= �ϑ �Z �v �� �;� �6� ��h  �|� ��3 � �t  �h8 郓  ��3 ��x �4�  �߈ �
  �e^  �0� �K� �6 �1 �� �w �� �� �� �s! ��^  ��� �|3 �� �O �5� ��c  �KP �V �q ��� �'� �2� �a �� �C� �� 驹 �4n  �_� ��7 酒 �o  �+T ��� �Q� �2 鷲 �3 ��  �}  �� �] �i �) �o� �z� �u� �0�  �5  �� �� ��� � 钺 �-�  �H� ��2 �� �~ ���  � ��� 饼  逿 �W4 �� �!� ��� �1 �2� �2 �� �� �� ��� �� 韙 �ڔ �5 �� �j �6�  �a �� �'�  �҂  �M �� �c �>� �Y�  �t�  �� �j� ��  适  �;�  �f� �a�  �� �8 �a �} �� ��� � �y�  �T7 �on �J� �> �pZ �{ �F� �1� 霛 �� ��� �m�  �� �Ӹ  �> �m  �t�  ��t 骵 饈 鐁  �[	 �ƾ ��2 �[ �m �� �] �ش ��> ��e ��  �4�  �0 �� �5U �0 �k& �N �A�  �2 �G �3 ��� � �ӧ �{ ��� �T� � �� ��i �:1 ��6 � ���  錴 �'_ �7 靜 ��� �S� �% �� �T\  � �- 酒 �  ��R �&�  ��  �L �; �"� �� 鸆 ��� 鞐  �y  �4Z  �/ �1 ��� ���  �� �M ��r �< ��j  ��^ �� ��V �C� 龔 �yW �Ĺ �� �J� �E� �~ �;� ��� ��	 �� ��� 钯 �� �(� �� �.  ��� �d�  �l  �z? �u& �  �۱  �&�  �Q�  �, �2 �r  �]/ �x� �C �.� ��  �� �l �j  �u � 3 �k�  �f� �1�  �̈  ��  �"� �m� �} �4 �~ �y� �Tp �?� �� �4 �- � �Ʈ  �� �\�  �w�  �b� �l �(� 飴 �  �) ��. �� �~ �e! �� � 閙 �qK �l� �'�  ���  �] �  ��  ���  �9 �d� �_  �z�  镜  �\  � 醏 �As ��� �w� �r� ���  �T �� �� ��  �tT �� �
 �� �0� �+ �� �!� �̰ �� �B{ 鍎  �H �c� �Nu  �Y �t� �o' �:� �� �- �;8 �6o  �� �s ���  �2 ��� �8� ��I �� � �t�  �ߕ �
�  ��X ��� �� ��, �� ��� �G �� ��  �8d  铣 �Ng  �S  �V, 鿗 �� �% � �� ��, �. ��� �M �B9 ��  �	 �s< ��� ��  ��A ��e  �Z+ ��  � � �[ �f; �Q �L�  �� �� �� �) �S2 �� ��1 �t� �/� ��1 �_ �@� � . �&�  �1 �; �� 邗  �M 騶 �s� � �� � �ϕ  ��� �� �@ �s  �� �q �� 駟 � ��]  ��s ��  �� �i� ��4 �y  ��( 酢  ��� �� �v �A� �,@ �� �� �=< �c 鳨 �~� �9� �dJ �/ �z0 �� ��_ �;S � �qs  �� �Gc ���  �}� �� �� �.Y ��K �4� �j �� �%7 �0�  �3* �f� ��� �l �'� �3 �� ��  �g ��4 �� � �?G ��l  �M* ��  �k�  ��  �m �<� �G� �u  ��) �h �# �> �i( �j � �: � �3 �k� �� ��u � �y �B� ���  �� � �� �� �� �� ��) ��? �@�  �{� �� �q� �* ��) �b� �-G �a ��}  �>{ ��  �4�  �/w �z� 镀 �p�  �� �~  �� �) ���  �* 魌 �X�  �m  � ��V ��  �|  �Z� 镉 �� 雌  ��( �� �l� ��B ���  �� �(� 鳄 ��M �i �� �_� �� 酿 �@ ��
 ��b �ѓ  ��  �� �R� �m ���  �> �.�  ��g �� �1 �� �u � q �K2 �6� ��0 �|: � �B8 �}u ��)  ��( �Ό �Yw �� �� �Z�  �;( �P� ��  �� �� �,� �' �B�  ��' �Hq �q  ��, ��8 �� �o� �j9 �u; �P�  �z  �1 � 鬽 �w �2� �=, �� �#� �� ��
 ��T �� �JW ��- � P  ��� �&�  �< ���  ��r  �� ��M � 飚 �^ ��, �:+ �ϵ �:
 � � � �k �6{  �' �<�  �'� �b�  ��N  �x- ��Y �. �p  �& �- 骔  �� �@R  �& �^  ��� �,� �W� �+ �b �x�  ��k �ދ �#& �t" �o- �� ��  ��] �[^  �v� �f �� ��J 邶  �� �o  �Cp �ޚ  ��& �T& �?� ��- �u �p� �{� �� �{% �� �8 鲭  �� �ؔ �S� �~� �	�  �< �[% �� �G �P�  �ˣ  �63 �a| �� 闋 �� �� �  �C� ��  �)% �> ���  骔 �- ��$ �G �F� �K �. ��  邹 �� �(� ��� �� �ym �4� �� ���  �u  �@| �+�  閷 �a� �|X �g& ��  �" �X �� �x ��5 �4� ��� �J7 �%�  ��� �u  �	 �^ � �w �R� �K �h% �� ��� �% ��B �/� �:� �5�  ���  �� �fj ��� �< �7N  ��s �$ �^ 郥  �l% �9� �T�  ��  ��\ �D �� �[� ��  � �� �@ �B) ��M �( �#� �>Y �i) �4� ��  �Z�  ��$ �� �� �&� �q� �N  闪 �"� �]�  ��W �< � �� ��  �� �*� 鵝 �p� �+� ��  �Q�  �l� �W �2� ��Y � �sq �2 �9� �t� �?�  �z�  �]  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������E���Ex��M�U;������EE�E��_^[���   ;��������]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�UR�EP�M������_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�UR�EP�M������_^[���   ;��#�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��(����6   ������Y�M��E�E�j�M��T����   _^[���   ;��v�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�BH���   �у�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ������9   ������Y�M��E�E�M������E�j h�  �M�����������$h�  �M�腹������<�$h�  �M��l�������<�$h�  �M��S�������<�$h�  �M��:����   _^[���   ;�������]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M��P0��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP�DX�Q�M��B,��;�����_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q@�B,�Ѓ�;�����_^[���   ;�������]����������������������������U����  SVWQ��(����6  ������Y�M��M�����E�E�E��M�������EԋM������EȋE�E��M������E��M��X����E�j h�  ��@���P�M�������������4�����@���������4��� ��  �M����������$�����$�����$��\�������P�����$�����$�����$��|����x���P�M����j�M�����M�蘽���M��?�����uǅ����    �M������������m  �E�P����������jj hgnlf������Q�U�R�����������������j hH=��h����O����E�P��h����)���P��P�������j j j �M��������������M��������������P���P�M���������������D����M�������������8����M������������M��������c���j ��8���P��D���Q�M��i������f����M��Z������!���h�   h�   h�   h�   �M��7������2�����P���Pj j �M�������������M������������M�����j��M�5���h�<� @��4Ph?]j`������������������� t#h�jj������Q�F�����������,����
ǅ,���    ��,�����,���h�<� @��5Ph?]j`�h����������������� t#h�jj������Q������������,����
ǅ,���    ��,����� ���h�<� @��6Ph?]j`������������������ t#h�jj������Q�|�����������,����
ǅ,���    ��,��������h�<� @��7Ph?]j`������������������ t#h�jj������Q������������,����
ǅ,���    ��,���������E��@�B����������E��@�1��������������$ۅ�������$ۅ�������$������������,������P�Q�P�Q�P�Q�P�Q�@�A�����$ۅ�������$�������D�����,���ۅ,������$�����茽����,��������P�Q�P�Q�P�Q�P�Q�@�A�����$�������8�����,���ۅ,������$�������D�����(���ۅ(������$��0���������,�����0��
�H�J�H�J�H�J�H�J�@�B�����$�������8�����,���ۅ,������$ۅ�������$��P���誼����,�����H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��p����\����� ������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������������ ��������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������û���� �����0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������u����� �����H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������'�����������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������ܺ������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��0���莺���������0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��P����@����������H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��p���������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������觹������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������Y����������0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�����������������H���P�Q�P�Q�P�Q�P�Q�@�Aǅ����    �M����������������������� u;ǅ����    ��P����Ю����h����Ů���M�轮���M��g����������  ǅ����    �������U��������������� u;ǅ����    ��P����q�����h����f����M��^����M������������W  ǅ����    �������4��������������� uj j�������D��������������� uJ������P豮����ǅ���    ��P���������h����ڭ���M��ҭ���M��|����������  ǅ����    ���������������������;�8�����   ǅ����    ���������������������;�D���}X������P������Q������R������P������Q����������������P������Q������R������P������荰����Y���j jj�����P�����Q�� ���R��,���P������Q�M�8���������P胭������,��� t��,�������������Q�b�����ǅ,���    �� ��� t�� ����� ����� ���Q�4�����ǅ ���    ����� t�������,�����,���Q������ǅ���    ����� t�������8�����8���Q�ة����ǅ���    j�M�}�������������������豼����uFǅD���    ������荳����P����Ы����h����ū���M�轫���M��g�����D����  �E�P��P�������jj hgnlf��P���Q������R�B�������P����G���j h�<��l�������������P��l����l���P��T��������j j j �������&������#����������������������T���P�������������� �����H����������������������<����������˹�����<���������蹹����蔾��j ��<���P��H���Q������藹����蔵��������腹�����L���h�   h�   h�   h�   �������_������Z�����T���Pj j �������B�����������������0�����衯���M�!���j��M�W���h�<� @�   Ph?]j`��������h�����h��� t#h�jj��h���Q�f�����h�����,����
ǅ,���    ��,�����0���h�<� @�   Ph?]j`膷������t�����t��� t#h�jj��t���Q�������t�����,����
ǅ,���    ��,�����$���h�<� @�   Ph?]j`������������������ t#h�jj������Q蘣����������,����
ǅ,���    ��,��������h�<� @�   Ph?]j`踶���������������� t#h�jj������Q�1�����������,����
ǅ,���    ��,���������E��@�\����� ����E��@ �K��������������$����������,���ۅ,������$�� �������(���ۅ(������$������������0�����
�H�J�H�J�H�J�H�J�@�B�����$����������,���ۅ,������$��H����� ����D
��(���ۅ(������$�������u�����0��������P�Q�P�Q�P�Q�P�Q�@�A�����$��<����������T��,���ۅ,������$��H����� ����T��(���ۅ(������$������������0�����0���P�Q�P�Q�P�Q�P�Q�@�A�����$��<����������T��,���ۅ,������$�� �������(���ۅ(������$�������x�����0�����H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������*�����$������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��8����߯����$��������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��X���葯����$�����0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��x����C�����$�����H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������誮������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�������\����������0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�����������������H���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$������������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��8����u�������������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��X����'����������0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��x����٬���������H���P�Q�P�Q�P�Q�P�Q�@�Aǅ����    ������輱�������������������� ugǅ����    ��T���蛢����l���萢��������腢���������,�����P����o�����h����d����M��\����M������������U  ǅ����    ����������������������� ugǅ����    ��T���������l������������������������衩����P���������h����١���M��ѡ���M��{�����������  ǅ����    ������觼�������������� uj j������距�������������� uv������P�$�����ǅ����    ��T����X�����l����M����������B���������������P����,�����h����!����M������M��è���������  ǅ����    �����������������8�����
9�������   ǅ����    �����������������D�����
9�����}X������P������Q������R������P������Q�������4���������P������Q������R������P�������Σ����S���j jj�����P�����Q��$���R��0���P������Q�M�y���������P�Ġ������0��� t��0���������������Q裝����ǅ0���    ��$��� t��$���������������Q�u�����ǅ$���    ����� t�����������������Q�G�����ǅ���    ����� t�����������������Q������ǅ���    j�M辩����T����@�����l����5����������*����������Ѧ����P���������h����	����M������M�諦���   R��P�(�c���XZ_^[���  ;�謱����]�    0����   ����   h���   P���   �����   �����   �����   �����   �l���   �T���   �����   �����   �r2 bmp2 objPointCount pnts countToString cm2 r bmp objPolygonCount plys polycountToString cm �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E�����E����X�E����X�E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��E��E��E�X�E��E�X�E�_^[��]� �����������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��������E�P�MQ�DX�B�H�у�;��ۨ���E�_^[���   ;��Ȩ����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��]�����EPj��MQ�U�R�DX�H�Q�҃�;��6����E�_^[���   ;��#�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;�譧��_^[���   ;�蝧����]����������������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M��,���P�M��k����E�_^[���   ;��/�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M��B<��;��Ҧ��_^[���   ;��¦����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M��BL��;��Q���_^[���   ;��A�����]� �����������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   ��Ѓ�;��{���_^[���   ;��k�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;�����_^[���   ;��������]� ����������������������������������U����   SVWQ������:   ������Y�M��M��m�����E�P�M�Q�DX�B@�H$�у�;�聤���E�P�M蟢���M�謒���ER��P��� ���XZ_^[���   ;��I�����]� �   �����   �bc ���������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H�Q<�҃�;�誣��_^[���   ;�蚣����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B��  �у�;�����_^[���   ;��
�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�Bd��H  �у�;�薢��_^[���   ;�膢����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Qd�Bh�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�Hd�Q$�҃�;�覡��_^[���   ;�薡����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R�DX�Hd���   �҃�$;�����_^[���   ;��������]�  ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�Bd���   �у�;�膠��_^[���   ;��v�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��G���_^[���   ;�������]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�HH���   �҃�;�裟��_^[���   ;�蓟����]� �������������������������������U����   SVWQ��4����3   ������Y�M�h�  �M�����_^[���   ;��.�����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�BH���   �у�;��ƞ��_^[���   ;�趞����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M�臑��_^[���   ;��L�����]���������������������������U����   SVWQ��4����3   ������Y�M�h�  �M��҈��_^[���   ;�������]�����������������������������U����   SVWQ��4����3   ������Y�M��DX���   ��M��Bt��;�菝��_^[���   ;�������]������������������������������U���|  SVWQ�������_   ������Y�M������$h�  ������P�M��������T����]荍�����I����E��E��X�����$h�  ������P�M辛���������]؍����������E��E��X�����$h�  ������P�M脛����������]ȍ������Պ���E��E��X�����$h�  ������P�M�J�����覗���]�������蛊���E��E��X 3�_^[��|  ;��A�����]� �����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP�DX�Q�M����   ��;�衛��_^[���   ;�葛����]� �����������������������������U���,  SVW�������K   ������h'  �Ά����P�M��
����M��9�����uǅ����   �M��C����������   j hh=�������\���j hX=������J���j ������P�����������������P�����Qh �j	�U�Rh�� �R�����������������胤�������轇��������貇���M�誇��������R��P�x����XZ_^[��,  ;��\�����]Ë�   �����   �path �������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�褤�������_^[���   ;�譙����]����������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVW��0����4   ������h�<jh?]j(�l�������8�����8��� t��8����&�����0����
ǅ0���    ��0���_^[���   ;��ؘ����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M�軒���E�� |=�E�_^[���   ;��g�����]����������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�������E�_^[���   ;��������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E�� �=�E�_^[���   ;�藗����]����������������������U����   SVWQ��4����3   ������Y�M��M�辁��_^[���   ;��C�����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�y������E�_^[���   ;�茖����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��s����E�� L>�E�_^[���   ;��'�����]����������������������U����   SVWQ��4����3   ������Y�M��M�蝋��_^[���   ;��ӕ����]������������������U����   SVWQ��4����3   ������Y�M��M�艆���E��t�E�P�Y������E�_^[���   ;��l�����]� ������������������������U����   SVWQ��4����3   ������Y�M�襉���M���E�_^[���   ;�������]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P�֔�����E��     _^[���   ;�覔����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVW��@����0   ������=@X t��EP�@X��;��ѓ��_^[���   ;��������]��������������������������������U���   SVW��������   ������j h�>�������˚��P�#������E��������~����}� u��  j h�>�����藚��P�E�P�@�����������������C��������� t�  j h�>�� ����Y���P�\������E썍 ��������M��}��j h�>��P����(���P��8�����~����8���Pj�M��u�����8���蠚����P������j h�>����������P��h����~����h���Pj�M��0�����h����[����������z��j������薍��������Pj�M�������������'���j h�>�������u���P�������*~��������Pj�M������������������������}� t1�E�P�������x����M�Q������Rj�M��>���������譙���+�E�P�������G���������Qj�M��U���������耙���M����R��P�x'����XZ_^[��   ;��Z�����]�   �'����   �'sc �����������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q�DX���   �H$�у�;������E�_^[���   ;��Џ����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q�DX���   �H0�у�;��C����E�_^[���   ;��0�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;�趎��_^[���   ;�覎����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P�M����   ��;��3���_^[���   ;��#�����]� �������������������������������U����   SVW��@����0   ������DX���   �@X�DXǀ�   ��w����u3���   _^[���   ;�融����]�����������������������������U����   SVW��@����0   ������_^[��]������������U���`  SVW�������X   ������E�������������  #�������  tZ������ tB������t�  �������  �u  ��  �PX�Rx����u3���  �   ��  �   ��  ��  �E�E��E�    �	�E���E�E��M�;�  �E��H�U�<� u��hd?�E��H�U��P�-�������th\?�E��H�U��P��������u1j hD?������荓��������P�0v�����������=y���   h<?�E��H�U��P��������u>�E��H�U���    j h$?�������.���������P��u������������x���8h?�E��H�U��P�d������u�E��H�U���    �    �  ������   �E�E��} u�s�E��x t�hj h�>������襒��������P�M��	�'x��P������R�����P��t����P�&u����������3x���������(x���������x��3��3�_^[��`  ;��������]���������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   ������EP�M������EP�M��N����E�P�M�̑���M��w���ER��P�/�{��XZ_^[���   ;��Љ����]Ë�   /����   /s ��������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@ƻ�E�@8W��E�@<H��E�@@���E�@D��E�@H���E�@L^��E�@P���E�@l:��E�@X���E�@\˶�E�@`��E�@d+��E�@T&��E�@hq��E�@p���E�@t0��E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������������U���h  SVW�������Z   ������j h�   ��\���P蛇����j �EP�MQ�UR�EP��\���Q�b������E �E�h�   ��\���P�MQ�URj��~����R��P�05�[u��XZ_^[��h  ;�褃����]Ë�   85\����   D5np ���������������������������������������������������������U����   SVW��@����0   ������EP�M���   Q�UR��s����_^[���   ;�������]���������������������U���  SVWQ��\����i   ������Y�M��,r���M���E��8 u��   �EP��l�����q��j hl?�����������P��������q��j j���l���Q������R������P��r����P������Q�@}����P�����R�0}����P�E����l��������؈�c���������u����������t����������t����������t���������o����l�����t����c�����t�E�P�o�����E�_^[�Ĥ  ;��������]� ��������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�z�����M���E�_^[���   ;�������]� �������������������U����   SVWQ��4����3   ������Y�M��E�P�n����_^[���   ;�迀����]�����������������������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U����   SVW��@����0   ������E�DX�DX� _^[��]�����������������������������U����   SVW��@����0   ������E�8 t��E�Q�DX�B��у�;��	���E�     _^[���   ;���~����]�������������������������������U����   SVW��@����0   �������hﾭޡDX�H��@  �҃�;��~��_^[���   ;��~����]������������������������������U����   SVW��@����0   ������} t!��EP�DX�Q��@  �Ѓ�;��~��_^[���   ;��	~����]������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;��}��_^[���   ;��}����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B��  �у�;��;}��_^[���   ;��+}����]��������������������������U����   SVW��@����0   ������DX�H��   ��;���|��_^[���   ;���|����]����������������������U����   SVW��@����0   ������} t�E�x��u�   �3�_^[��]��������������������U����   SVW��<����1   ������=DX tE�}sǅ<���   �	�E��<�����j j ��<���Q�DX�B���   �у�;���{���j�EP�I   ��_^[���   ;���{����]���������������������������������������������������U����   SVW��4����3   ������}s�E   �E��P� o�����E��}� u3��:�} t�E��Pj �M�Q�l�����E�� �����E����E��HX   �E�_^[���   ;��{����]��������������������������������������������U����   SVW��<����1   ������=DX tE�}sǅ<���   �	�E��<�����j j ��<���Q�DX�B���   �у�;��tz���j�EP�������_^[���   ;��Tz����]���������������������������������������������������U����   SVW��<����1   ������=DX tE�}sǅ<���   �	�E��<�����j j ��<���Q�DX�B���   �у�;��y���j�EP�	�����_^[���   ;��y����]���������������������������������������������������U����   SVW��<����1   ������=DX tE�}sǅ<���   �	�E��<�����j j ��<���Q�DX�B���   �у�;���x���j�EP�I�����_^[���   ;���x����]���������������������������������������������������U����   SVW��4����3   ������} tF�E�E��=HX t�E�x��u�E��P�M��������E�P�DX�Q��Ѓ�;��4x��_^[���   ;��$x����]�����������������������������������U����   SVW��4����3   ������} tF�E�E��=HX t�E�x��u�E��P譀�������E�P�DX�Q��Ѓ�;��w��_^[���   ;��w����]�����������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;��#w��_^[���   ;��w����]����������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;��v��_^[���   ;��v����]����������������������������������U����   SVW��<����1   ������=DX tI�}sǅ<���   �	�E��<�����MQ�UR��<���P�DX�Q���   �Ѓ�;��v���j�EP�e�����_^[���   ;���u����]�����������������������������������������������U����   SVW��<����1   ������=DX ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P�DX�Q���   �Ѓ�;��Fu���[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P�DX�Q���  �Ѓ�;���t����EP�MQ�N�����_^[���   ;���t����]������������������������������������������������������������������������U����   SVW��0����4   ������} w�E   �=DX t0��EP�MQ�UR�DX�H���   �҃�;��2t����0����j�EP��������0�����0����M��E���thp?�t@��
P��a�����E�_^[���   ;���s����]�����������������������������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B��0  �у�;��[s��_^[���   ;��Ks����]��������������������������U����   SVW��0����4   ������} w�E   �=DX to�} t0��EP�MQ�UR�DX�H���   �҃�;���r����0����.��EP�MQ�UR�DX�H���  �҃�;��r����0�����0����E��j�EP��������E��E���thp?�x@��P�5`�����E�_^[���   ;��Ir����]������������������������������������������������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;���q��_^[���   ;��q����]����������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;��Sq��_^[���   ;��Cq����]����������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;���p��_^[���   ;���p����]����������������������������������U����   SVW��@����0   �������EP�DX�Q��Ѓ�;��sp��_^[���   ;��cp����]����������������������������������U����   SVW��@����0   ������DX�H���   ��;��p��_^[���   ;���o����]����������������������U����   SVW��@����0   �������E�Q�DX�B���   �у�;��o���E�     _^[���   ;��o����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q���   �Ѓ�;��o��_^[���   ;��
o����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B���   �у�;��n��_^[���   ;��n����]� ����������������������������������U����   SVW��@����0   ������DX�H����;��;n��_^[���   ;��+n����]��������������������������U����   SVW��@����0   �������E�Q�DX�B�H�у�;���m���E�     _^[���   ;��m����]��������������������������������������U����   SVW��@����0   �������E�Q�DX�B�H�у�;��Pm���E�     _^[���   ;��7m����]��������������������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q�DX�B���   �у�;��l�����x��������� ����t�������_^[���   ;��l����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   �B8�Ѓ�;��l��_^[���   ;��
l����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��k��_^[���   ;��k����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�H\�у�;��9k��_^[���   ;��)k����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H���   �҃�;��j��_^[���   ;��j����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B�HX�у�;��j��_^[���   ;��j����]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B �Ѓ�;��i��_^[���   ;��i����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B���   �у�;��*i��_^[���   ;��i����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q�B�Ѓ�;��h��_^[���   ;��h����]� �����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�DX�B��   �у�;��h��_^[���   ;��h����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M��B$��;��g��_^[���   ;��g����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M���x  ��;��&g��_^[���   ;��g����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M���|  ��;��f��_^[���   ;��f����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B�H(�у�;��-f��_^[���   ;��f����]� �������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�DX�Q�B`�Ѓ�(;��e��_^[���   ;��e����]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B�H,�у�;��e��_^[���   ;���d����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M���m����P�M��)M����Pj j �E�P�DX�Q�B4�Ѓ� ;��ud��_^[���   ;��ed����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;���c��_^[���   ;���c����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��c��_^[���   ;��}c����]����������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q�DX�B�H4�у� ;��c��_^[���   ;���b����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H�Q@�҃�;��b��_^[���   ;��vb����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�HD�у�;��	b��_^[���   ;���a����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�BL�Ѓ�;��a��_^[���   ;��}a����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�BL�Ѓ�;��a��_^[���   ;��a����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�BP�Ѓ�;��`��_^[���   ;��`����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�HT�у�;��9`��_^[���   ;��)`����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�HT�у�;��_��_^[���   ;��_����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H���   �҃�;��3_��_^[���   ;��#_����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P�DX�Q���   �Ѓ�;��^��P�M��^���� ����f���E_^[���   ;��^����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q�DX���   �H�у�;��^���E�_^[���   ;���]����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�Bh�Ѓ�;��}]��_^[���   ;��m]����]����������������������������U����   SVW��0����4   ������h�?�|@��Ph?]h�   �bc������8�����8��� t��8����dg����0����
ǅ0���    ��0���_^[���   ;���\����]���������������������������������������������U����   SVW��$����7   ������E�8 t?�E���8�����8�����,�����,��� tj��,����je����$����
ǅ$���    �E�     _^[���   ;�� \����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��M��tP���E��t�E�P�M�����E�_^[���   ;��[����]� ������������������������U����   SVWQ��4����3   ������Y�M��M����2V���M���^���E�_^[���   ;��5[����]��������������������U����   SVWQ��(����6   ������Y�M��M��a���E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��Z����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M���T���M����~R��_^[���   ;��HZ����]�����������������������U����   SVWQ��4����3   ������Y�M��M���L��_^[���   ;���Y����]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E����Xp�E��@x�����E��@|   _^[��]������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	�p^���E��     �E��x` t�E���`P��F����_^[���   ;���X����]������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 th�?��@��P�FF�����E��x` th�?��@��P�'F�����M��R���M���[���E�P�M���dQ�U��BxP�MQ�U���`R�_�����M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�E�����E��@|�   �E��xd ��   �E���pP�M���hQ�UR�V������u(�E��@h    �E����Xph�?��@��P�JE�����EP�M����_��j j j�E���P�M��	�\���U��B|�E��x|t�M��Q���E��@|��E��@x�����E��@|_^[���   ;��W����]� ������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M���P���M���Y��_^[���   ;��KV����]��������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	�-[���U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;��mU����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap��E��xd t�E��@h��E��x|u�   �3�_^[��]� ��������������������������������U����   SVW��@����0   ������DX�H����;��{T��_^[���   ;��kT����]��������������������������U����   SVW��@����0   �������E�Q�DX�B�H�у�;��T���E�     _^[���   ;���S����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q�DX�B�H�у� ;��qS��_^[���   ;��aS����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�H�у�;���R��_^[���   ;���R����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��}R��_^[���   ;��mR����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H�Q�҃�;��R��_^[���   ;���Q����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��<�����M��<���H �G@��;��|Q��_^[���   ;��lQ����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M���;�����M���;���H �GD��;���P��_^[���   ;���P����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M��z;���xH u3��#�M��h;�����M��^;�����H �FH��;��VP��_^[���   ;��FP����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M���:���xL u3��/��EP�MQ�UR�M���:�����M���:���H �GL��;��O��_^[���   ;��O����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M��J:���xP u����3��EP�MQ�UR�EP�M��%:�����M��:���H �WP��;��O��_^[���   ;��O����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M��9���xT u����+��EP�MQ�M��9�����M��9���H �WT��;��}N��_^[���   ;��mN����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��M��
9���xX u����'��EP�M���8�����M���8���H �WX��;���M��_^[���   ;���M����]� �����������������������������U���  SVWQ�������C   ������Y�M��} t<�M��G8����E�P�M��f8�����M��\8���H �WL��;��VM���M��M��;���} t?��������Q��P�M�v=���������K:���M��8���@@�EЃ}� t�E�P�M�K=��R��P��k�>��XZ_^[��  ;���L����]� �I    �k����   lbc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�DX�B�H�у�;��9L���E�_^[���   ;��&L����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q�B�Ѓ�;��K���E�_^[���   ;��K����]�������������������������U����   SVWQ��4����3   ������Y�M��M��Z6���x` u� }  �'��EP�M��?6�����M��56���H �W`��;��/K��_^[���   ;��K����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��5�����M��5���H �WH��;��J��_^[���   ;��J����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�j�EP��R���������P�M��9���E�M�2��;E��M�DS��;E�~������3��EP�MQ�UR�EP�M���4�����M���4���H �WD��;���I��_^[���   ;���I����]� ���������������������������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M��4���xP u������;��EP�MQ�UR�EP�MQ�UR�M���3�����M���3���H �GP��;���H��_^[���   ;���H����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��j3���xT u������+��EP�MQ�M��K3�����M��A3���H �WT��;��;H��_^[���   ;��+H����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M���2���xX u�'��EP�M��2�����M��2���H �WX��;��G��_^[���   ;��G����]� ��������������������������������U����   SVW�� ����8   ������M�� D���E�P�MQ�R������t�}� u3���E�P�M�Q�U�R�E�P�M��J��R��P��q�8��XZ_^[���   ;���F����]ÍI    �q����   �qdat ����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVWQ������<   ������Y�M��M�S0���M��=����uh�?��@��P�3����3��   �E�    ��E�P�M�Q�UR�E�P�DX�Q���   �Ѓ�;��E����u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�)3���͍E�P�>�����   R��P��s��6��XZ_^[���   ;��E����]�    �s����   �s����   �sarr count ����������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M��4���M��;����uh�?��@��P�2����3��   �E�    ��E�P�M�Q�UR�E�P�DX�Q���   �Ѓ�;��D����u3��i�}� u3��_�E�    �	�Eԃ��EԋE�;E�}4�EԋM��<� t�EԋM���� ;����u�ϋEԋM���R�M�[J��뻍E�P��<�����   R��P�`u�+5��XZ_^[���   ;��tC����]�    hu����   �u����   �uarr count ��������������������������������������������������������������������������������������U����   SVW��@����0   ������DX�H��   ��;��B��_^[���   ;��B����]����������������������U����   SVW��@����0   �������E�Q�DX�B��$  �у�;��MB���E�     _^[���   ;��4B����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�DX�B��(  �у�;���A���E�_^[���   ;��A����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�DX�B��,  �у�;��FA��_^[���   ;��6A����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�DX�B��,  �у�;���@�������_^[���   ;��@����]� ���������������������������U����   SVW��@����0   ������DX�H��0  ��;��W@��_^[���   ;��G@����]����������������������U����   SVW��@����0   ������DX�H��4  ��;���?��_^[���   ;���?����]����������������������U����   SVW��@����0   ������DX�H��p  ��;��?��_^[���   ;��?����]����������������������U����   SVW��@����0   ������DX�H��t  ��;��7?��_^[���   ;��'?����]����������������������U����   SVWQ��0����4   ������Y�M��} t�M�J;����0����
ǅ0���    ��0���P�M�Q�DX�B��8  �у�;��>��_^[���   ;��>����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��<  �у�;���=��_^[���   ;���=����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q��@  �Ѓ�;��N=��_^[���   ;��>=����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H��D  �҃�;���<��_^[���   ;���<����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��H  �у�;��V<��_^[���   ;��F<����]� ����������������������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R�DX�H��L  �҃�;���;��P�M�C���� �����(���E_^[���   ;��;����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q��T  �Ѓ�;��:;��_^[���   ;��*;����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��l  �у�;���:��_^[���   ;��:����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q��P  �Ѓ�;��J:��_^[���   ;��::����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��X  �у�;���9��_^[���   ;���9����]� ����������������������������������U����   SVW��@����0   ������DX�H��\  ��;��g9��_^[���   ;��W9����]����������������������U����   SVW��@����0   �������E�Q�DX�B��`  �у�;���8���E�     _^[���   ;���8����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H��d  �҃�;��g8��_^[���   ;��W8����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H��h  �҃�;���7��_^[���   ;���7����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��g+��_^[���   ;��_7����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��7����]������������������U����   SVWQ��4����3   ������Y�M��EP�M��*��_^[���   ;��6����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��S6����]������������������U����   SVW��4����3   ������j�[   ���E��}� t	�E��x u3���E���H��;���5��_^[���   ;���5����]������������������������������U����   SVW��@����0   ������hLX�EPh.D �� ����_^[���   ;��z5����]�������������������������U����   SVW��4����3   ������j�{������E��}� t	�E��x u���EP�M��Q�҃�;��
5��_^[���   ;���4����]�����������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u���� ��EP�MQ�UR�E�M��P��;��*4��_^[���   ;��4����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u������EP�U�M��B��;��3��_^[���   ;��3����]� ������������������������������U����   SVWQ��(����6   ������Y�M�j�v������E�}� t	�E�x u������EP�MQ�U�M��B��;���2��_^[���   ;���2����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u���� ��EP�MQ�UR�E�M��P��;��Z2��_^[���   ;��J2����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j �6������E�}� t	�E�x  u���E�M��P ��;���1��_^[���   ;��1����]����������������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u���EP�MQ�U�M��B$��;��11��_^[���   ;��!1����]� �����������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u������E�M����   ��;��0��_^[���   ;��0����]��������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u������E�M����   ��;���/��_^[���   ;���/����]��������������������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3����E�M��P(��;��g/��_^[���   ;��W/����]��������������������������������������U����   SVWQ��(����6   ������Y�M�j,�F������E�}� t	�E�x, u���E�M��P,��;���.��_^[���   ;���.����]����������������������������������������U����   SVWQ��(����6   ������Y�M�j0�������E�}� t	�E�x0 u���E�M��P0��;��I.��_^[���   ;��9.����]����������������������������������������U����   SVWQ��(����6   ������Y�M�j4�&������E�}� t	�E�x4 u���EP�MQ�U�M��B4��;��-��_^[���   ;��-����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u���EP�MQ�U�M��B8��;��!-��_^[���   ;��-����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j<�������E�}� t	�E�x< u�$��EP�MQ�UR�EP�U�M��B<��;��,��_^[���   ;��y,����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�j@�f������E�}� t	�E�x@ u���EP�MQ�U�M��B@��;���+��_^[���   ;���+����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jD��������E�}� t	�E�xD u�$��EP�MQ�UR�EP�U�M��BD��;��Y+��_^[���   ;��I+����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�jH�6������E�}� t	�E�xH u���EP�MQ�U�M��BH��;���*��_^[���   ;��*����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jL�������E�}� t	�E�xL u���EP�MQ�U�M��BL��;��1*��_^[���   ;��!*����]� �����������������������������U����   SVWQ��(����6   ������Y�M�jP�������E�}� t	�E�xP u�$��EP�MQ�UR�EP�U�M��BP��;��)��_^[���   ;��)����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�jT�v������E�}� t	�E�xT u�$��EP�MQ�UR�EP�U�M��BT��;���(��_^[���   ;���(����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�jX��������E�}� t	�E�xX u�(��EP�MQ�UR�EP�MQ�U�M��BX��;��U(��_^[���   ;��E(����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j\�6������E�}� t	�E�x\ u�(��EP�MQ�UR�EP�MQ�U�M��B\��;��'��_^[���   ;��'����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j`�������E�}� t	�E�x` u�$��EP�MQ�UR�EP�U�M��B`��;��'��_^[���   ;��	'����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�jd��������E�}� t	�E�xd u�$��EP�MQ�UR�EP�U�M��Bd��;��y&��_^[���   ;��i&����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�jh�V������E�}� t	�E�xh u�,��EP�MQ�UR�EP�MQ�UR�E�M��Ph��;���%��_^[���   ;���%����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�jl�������E�}� t	�E�xl u�,��EP�MQ�UR�EP�MQ�UR�E�M��Pl��;��!%��_^[���   ;��%����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�jp��������E�}� t	�E�xp u� ��EP�MQ�UR�E�M��Pp��;��}$��_^[���   ;��m$����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M�jt�V������E�}� t	�E�xt u3����EP�U�M��Bt��;���#��_^[���   ;���#����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jx��������E�}� t	�E�xx u3����E�M��Px��;��W#��_^[���   ;��G#����]��������������������������������������U����   SVWQ��(����6   ������Y�M�j|�6������E�}� t	�E�x| u3����E�M��P|��;���"��_^[���   ;��"����]��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u�7��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�M����   ��;��"��_^[���   ;�� "����]�  ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u�'��EP�MQ�UR�EP�U�M����   ��;��`!��_^[���   ;��P!����]� ��������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u�#��EP�MQ�UR�E�M����   ��;�� ��_^[���   ;�� ����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;�� ��_^[���   ;�� ����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��'��EP�MQ�UR�EP�U�M����   ��;��n��_^[���   ;��^����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u3��$����E�$�EP�U�M����   ��;�����_^[���   ;������]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u�����EP�U�M����   ��;����_^[���   ;��
����]� ��������������������������������������U����   SVW��4����3   ������h�   ��������E��}� t-�E����    t!��EP�MQ�U����   �Ѓ�;�����3�_^[���   ;��k����]������������������������������������������U����   SVW��4����3   ������h�   �X������E��}� t1�E����    t%��EP�MQ�UR�E����   �у�;������3�_^[���   ;�������]��������������������������������������U����   SVW��4����3   ������h�   �������E��}� t6�E����    t*����E�$�EP�MQ�U����   �Ѓ�;��6���3�_^[���   ;��"����]���������������������������������U����   SVW��4����3   ������h�   �������E��}� t1�E����    t%��EP�MQ�UR�E����   �у�;�����3�_^[���   ;������]��������������������������������������U����   SVW��4����3   ������h�   �x������E��}� t/�E����    t#��EP�MQ�UR�E����   �у�;�����3�_^[���   ;�������]����������������������������������������U����   SVW��4����3   ������h�   ��������E��}� t-�E����    t!��EP�MQ�U����   �Ѓ�;��_����M�|%��_^[���   ;��E����]������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B8�HD�у�;��i��_^[���   ;��Y����]� �������������������������������������U����   SVW��@����0   ������DX�H8��Q<��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������E�Q�DX�B8�H@�у�;�����E�     _^[���   ;��w����]��������������������������������������U����   SVW��@����0   ������DX�H8����;����_^[���   ;������]��������������������������U����   SVW��@����0   �������E�Q�DX�B8�H�у�;�����E�     _^[���   ;������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q8�B�Ѓ�;��!��_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H8�Q�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q8�B�Ѓ�;��-��_^[���   ;������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B8�H �у�;����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H8�Q$�҃�;��*��_^[���   ;������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P�DX�Q8�B�Ѓ�;����_^[���   ;������]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H8�Q(�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q8�B,�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q8�B�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�DX�H8�Q�҃�;����_^[���   ;��z����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H8�Q0�҃�;����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q8�B4�Ѓ�;����_^[���   ;��q����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B8�H8�у�;��	��_^[���   ;�������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q��x  �Ѓ�;����_^[���   ;��s����]����������������������������������U����   SVW��@����0   �������EP�MQ�DX�B��|  �у�;����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;��+��_^[���   ;������]��������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP�DX�Q�B,�Ѓ�;��R��_^[���   ;��B����]���������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP�DX�Q���  �Ѓ�;�����_^[���   ;������]��������������������������������������U����   SVW��(����6   ������M�������E�P�DX�Q�B8�Ѓ�;��J���E�P�M����M��]����ER��P��������XZ_^[���   ;������]�   ȫ����   ԫstr ����������������������������������������U����   SVW��@����0   ������DX�H��Q<��;����_^[���   ;������]�������������������������U����   SVW��@����0   �������EP�MQ�DX�B�H@�у�;��.��_^[���   ;������]�����������������������������U����   SVW��@����0   ������DX�H��QD��;�����_^[���   ;������]�������������������������U����   SVW��@����0   ������DX�H��QH��;��j��_^[���   ;��Z����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H�QL�҃�;���
��_^[���   ;���
����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B�HP�у�;��
��_^[���   ;��~
����]�����������������������������U����   SVW��@����0   �������EP�DX�Q��<  �Ѓ�;��
��_^[���   ;��
����]������������������������������U����   SVW��@����0   �������EP�DX�Q��,  �Ѓ�;��	��_^[���   ;��	����]������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP�DX�Q���   �Ѓ�;��	��_^[���   ;��	����]���������������������������������������U����   SVW��@����0   ������DX�H�􋑼   ��;����_^[���   ;������]����������������������U����   SVW��@����0   ������DX�H���  ��;��G��_^[���   ;��7����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�2  �DX�B���   �у�;�����_^[���   ;������]�����������������������������������������U����   SVW��@����0   �������EP�DX�Q�B�Ѓ�;��R��_^[���   ;��B����]���������������������������������U����   SVW��@����0   �������EP�DX�Q��\  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������<   ������EPj h@���������P�M�Q�"����������������E�P�DX�Q�B�Ѓ�;��D���M��c���R��P��������XZ_^[���   ;������]Ð   ������   ̲s ��������������������������������������������������U����   SVW��@����0   �������EP�DX�Q�BT�Ѓ�;����_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP�DX�Q�BX�Ѓ�;��"��_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP�DX�Q�B\�Ѓ�;����_^[���   ;������]���������������������������������U����   SVW��@����0   ������DX�H��Q`��;��J��_^[���   ;��:����]�������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   ������DX�H��Qd��;��z��_^[���   ;��j����]�������������������������U����   SVW��@����0   ������DX�H��Qh��;����_^[���   ;��
����]�������������������������U����   SVW��@����0   �������EP�DX�Q�Bl�Ѓ�;����_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP�DX�Q�Bp�Ѓ�;��B��_^[���   ;��2����]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H�Qt�҃�;�����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP�DX�Q��D  �Ѓ�;��_��_^[���   ;��O����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q��  �Ѓ�;��� ��_^[���   ;��� ����]����������������������������������U����   SVW��@����0   �������EP�MQ�DX�B�Hx�у�;��n ��_^[���   ;��^ ����]�����������������������������U����   SVW��@����0   �������EP�MQ�DX�B��@  �у�;������_^[���   ;��������]��������������������������U����   SVW������9   ������M�������E�P�MQ�DX�B�H|�у�;������E�P�M����M��W����ER��P�������XZ_^[���   ;��N�����]�   ������   ��fn �����������������������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B���   �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B��h  �у�;��K���_^[���   ;��;�����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q��d  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��X���_^[���   ;��H�����]�����������������������U����   SVW��@����0   ������DX�H�􋑄   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ�DX�B��l  �у�;�����_^[���   ;��{�����]��������������������������U����   SVW��@����0   �������EP�DX�Q��   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��$����7   ������M��"�����E�P�DX�Q���   �Ѓ�;��7����E�P�M�U����M��b����ER��P�Խ����XZ_^[���   ;��������]Ð   ܽ����   �bc �����������������������������������������������������U����   SVW��@����0   ������DX�H��`  ��;��w���_^[���   ;��g�����]����������������������U����   SVW��@����0   �������EP�DX�Q��  �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVW�� ����8   �������EP��$���Q�DX�B���   �у�;������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��`�����]�����������������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ�DX�B���   �у�;��i���_^[���   ;��Y�����]����������������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���   �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���   �҃�;��x���_^[���   ;��h�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��(���_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���   �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�DX�B���   �у�;��K���_^[���   ;��;�����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B���   �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�DX�Q���   �Ѓ�;��o���_^[���   ;��_�����]������������������������������U����   SVW��@����0   �������EP�DX�Q���   �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�DX�Q���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�DX�Q���   �Ѓ�;�������u3���E�R��P�������XZ_^[���   ;��������]�   ������   (�����   !�����   �data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�DX�Q���   �Ѓ�;�������u3���E�R��P�������XZ_^[���   ;��������]�   ������   �����   �����   �data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�DX�Q���   �Ѓ�;��.�����u3���E�R��P�������XZ_^[���   ;�������]�   ������   �����   �����   ��data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP�DX�Q��8  �Ѓ�;��O���_^[���   ;��?�����]������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�>���P�U�R�DX�H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M����P�U�R�DX�H0���   �҃�(;�����_^[���   ;��������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�DX�Q0���   �Ѓ�(;�����_^[���   ;�������]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B0���   �у�;�����_^[���   ;��z�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q0���   �Ѓ�;��
���_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H0���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�DX�B0���   �у�;��
���_^[���   ;��������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q0���   �Ѓ�;�����_^[���   ;��z�����]�������������������������U����   SVW��@����0   ������DX�H0�􋑤   ��;��'���_^[���   ;�������]����������������������U����   SVW��@����0   �������E�Q�DX�B0���   �у�;������E�     _^[���   ;�������]�����������������������������������U����   SVW��@����0   �������EP�DX�Q��H  �Ѓ�;��?���_^[���   ;��/�����]������������������������������U����   SVW��@����0   �������EP�DX�Q��T  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   ������DX�H��p  ��;��g���_^[���   ;��W�����]����������������������U����   SVW��@����0   ������DX�H���  ��;�����_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;��/���_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q���  �Ѓ�;��C���_^[���   ;��3�����]����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�DX�B���  �у�;�����_^[���   ;�������]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P�DX�Q��X  �Ѓ�;��@���P�M�i�����,����)����E_^[���   ;�������]����������������������������������������U����   SVW������=   ������j hLGOg���������PhicMC�E�P�.����������������M��U�����u�M�W����M������E��M��4���P�M�����M��d����ER��P��������XZ_^[���   ;��C�����]Ð   ������   ��dat ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   �BT�Ѓ�;�����_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ�DX�B��  �у�;��;���_^[���   ;��+�����]��������������������������U����   SVW��@����0   �������EP�DX�Q��\  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW������9   ������EP��MQ�� ���R�DX�H��t  �҃�;��U������>����� ����(����E_^[���   ;��0�����]�������������������������������U����   SVW��(����6   �������EP��,���Q�DX�B���  �у�;������P�M������,���������E_^[���   ;�������]��������������������������������U����   SVW��(����6   �������EP��,���Q�DX�B���  �у�;��8���P�M�������,����K����E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;��?���_^[���   ;��/�����]������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ�DX�B���  �у� ;��C���_^[���   ;��3�����]����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�DX�H���  �҃�$;�����_^[���   ;�������]�������������������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q�DX�B��t  �у�;��*���P�M�������,����=����E_^[���   ;�������]����������������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q�DX�B���  �у�;�����P�M������,����u����E_^[���   ;��e�����]������������������������������������U����   SVW��@����0   �������EP�DX�Q��8  �Ѓ�;������_^[���   ;��������]������������������������������U����  SVW��(����6  �����󫡐A3ŉE��E�E�E�P�MQh   ������R�������������Ph@�DX�Q��4  �Ѓ�;��[����E�    R��P��������XZ_^[�M�3��[������  ;��)�����]ÍI    ������   ��t ��������������������������������������������������������������U����   SVW��4����3   ������} 3��^�EP�MQ�UR�EP�D������E��}� |�E��9E�|/�}� }h @��@��P�7������EE�@� �E���E��E�_^[���   ;��8�����]���������������������������������������U����   SVW��(����6   �������,���P�DX�Q��  �Ѓ�;������P�M������,���������E_^[���   ;�������]������������������������������������U����   SVW��(����6   �������,���P�DX�Q��  �Ѓ�;��<���P�M������,����O����E_^[���   ;�������]������������������������������������U����   SVW������=   �������"�����u�\h���M������EPh���M�� ����EPh���M������j �E�PhicMC�����Q�������������n����M�����R��P��������XZ_^[���   ;��H�����]Ë�   ������   ��msg ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M��P4��;�����_^[���   ;�������]� �������������������������������������U����   SVW������=   ������������u�M������E�^h!���M������EPh!���M��u���j �E�PhicMC�����Q�������������P�M����������������M������ER��P���r���XZ_^[���   ;�������]Ð    �����   ,�msg ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   �BH�Ѓ�;�����_^[���   ;��
�����]�������������������������U����   SVW������=   �������"�����u�M�Q����E�^h����M������EPh����M������j �E�PhicMC�����Q���������o���P�M�B���������d����M������ER��P��������XZ_^[���   ;��;�����]Ð   ������   ��msg ����������������������������������������������������������������U���   SVW�� ����@   ������������u3��^h#���M������EPh#���M������j �E�PhicMC�����Q�������������������������`����M����������R��P��������XZ_^[��   ;��4�����]Ë�   ������   ��msg ��������������������������������������������������������U���   SVW�� ����@   ������������u3��^hs���M������EPhs���M������j �E�PhicMC�����Q�������������������������`����M����������R��P��������XZ_^[��   ;��4�����]Ë�   ������   ��msg ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;��|�����]���������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��@  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   ������E�8 t#��E�Q�DX�B��D  �у�;��%����E�     _^[���   ;�������]���������������������������U����   SVW��@����0   �������EP�DX�Q��H  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�DX�Q��L  �Ѓ�;��?���_^[���   ;��/�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��P  �҃�;������_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��T  �҃�;��X���_^[���   ;��H�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��X  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��\  �҃�;��x���_^[���   ;��h�����]�����������������������U����   SVW��@����0   ������DX�H��d  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP�DX�Q��h  �Ѓ�;�����_^[���   ;�������]��������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B��l  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   ������DX�H�􋑄  ��;�����_^[���   ;�������]����������������������U����   SVW��$����7   �������EP��(���Q�DX�B���  �у�;��H���P�M�i�����(����s����E_^[���   ;��!�����]��������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;��O���_^[���   ;��?�����]������������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;��o���_^[���   ;��_�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;��x�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��l  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;��?���_^[���   ;��/�����]������������������������������U����   SVW��@����0   �������EP�MQ�DX�B��$  �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�DX�Q��(  �Ѓ�;��_���_^[���   ;��O�����]������������������������������U����   SVW��@����0   �������EP�DX�Q��,  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   ������DX�H��0  ��;�����_^[���   ;��w�����]����������������������U����   SVW��@����0   ������DX�H��<  ��;��'���_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   ������DX�H���  ��;��G���_^[���   ;��7�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��4����3   ������j �M�����E��}� t�E�P�<������E�P�ɿ����R��P��������XZ_^[���   ;��D�����]Ë�   ������   ��c ������������������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ�DX�B��  �у� ;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   ������DX�H��P  ��;��7���_^[���   ;��'�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��`  �҃�;������_^[���   ;�������]�����������������������U����   SVWQ��4����3   ������Y�M��E���P�������_^[���   ;��\�����]���������������������������U����   SVW��@����0   �������EP�DX���   ���   �Ѓ�;������_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M���j j��DX�P�M��B��;������E�_^[���   ;��{�����]��������������������������U����   SVWQ��4����3   ������Y�M���j �EP�DX�Q�M��B��;������E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EPj��DX�Q�M��B��;������E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M��Z���_^[���   ;��#�����]������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M觹���E�_^[���   ;��������]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P�M����   ��;��c���_^[���   ;��S�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�H�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B�H�у�;��i��������_^[���   ;��R�����]� ������������������������������U����   SVWQ��(����6   ������Y�M��EP�M������E�M��1���_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   �BX�Ѓ�;��z���_^[���   ;��j�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bt��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M�����_^[���   ;�薾����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P�M��Bl��;��&���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M������_^[���   ;�覽����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��c����E�EP�M�賩��_^[���   ;��0�����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX���   �H`�у�;��Ƽ��_^[���   ;�趼����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��J���_^[���   ;��:�����]� ����������������������U����   SVWQ��(����6   ������Y�M���EP�DX�Q�M����   ��;��ڻ���E�}� u3���M��^���_^[���   ;�赻����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX���   �B�Ѓ�;��J���_^[���   ;��:�����]�������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����  SVW������z   ������M�?�����tj �EP�MQ誣������u3��Sj h   ������P蕽�����EP�M Q�UR�EP������Q�   ��h   ������P�MQ�URj�Դ����R��P�,��]���XZ_^[���  ;�覹����]�   4�����   @�np �������������������������������������������������������������U����   SVW��@����0   ������j �EP�MQ�UR�EP�MQ�������Eǀ�   ���Eǀ�   ��Eǀ�   ��_^[���   ;��۸����]�����������������������������������������̋�`L����������̋�`D����������̋�`H�����������U����   SVW��<����1   ������} t�E��<�����PX�G�����<�����<���Q�UR�EP襱����_^[���   ;�������]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��_���_^[���   ;�������]������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q�DX�B<�H�у�;�蕶���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� �������������
ǅ���    �E��@    _^[���   ;�� �����]���������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�蘨���E��t�E�P�y������E�_^[���   ;�茵����]� ������������������������U����   SVWQ������?   ������Y�M������P賥����P�M������������������������_^[���   ;�������]���������������������������U����   SVWQ��$����7   ������Y�M��E��x ufhp@��@��Ph?]j���������,�����,��� t�MQ��,���觼����$����
ǅ$���    �U���$����B�E��x u3��Q�E��x t�E�3Ƀ8 �����9��EP�DX�Q<��Ѓ�;��'����M���E��@   �E�3Ƀ8 ����_^[���   ;��������]� �����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@   �DX�H<��Q��;��k����M���E�3Ƀ8 ����_^[���   ;��I�����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �4�E��x u3��'��E��HQ�U��P�DX�Q<�B�Ѓ�;�跲��_^[���   ;�觲����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u�DX�H��#��EP�M��R�DX�H<�Q�҃�;��$���_^[���   ;�������]� ��������������������������������U����   SVW��@����0   ������PX����_^[���   ;�趱����]���������������������U����   SVW��@����0   ������EP�PX�n���_^[���   ;��b�����]�����������������U���  SVW�������B   ������EP�PX����P�M�����j h�@������d���j �E�P�����Q�M���������������������������������t�M�Y����M������E�9j�E�P�M��ɧ��j�j��EP�M�Q�M�������E�P�M�\����M�諝���ER��P�t����XZ_^[��  ;��`�����]Ë�   |����   �����   �str pos ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P�M��B@��;�薯��_^[���   ;�膯����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M��PH��;�����_^[���   ;��	�����]� �������������������������������������U���,  SVW�������K   ������EP�PX讙��P�M��y���j h�@�����������j �E�P������Q�M�覲�������������������葛����������t�M�����M��v����E�   j�E�P�M��V���j�j��EP�M�Q�M��N���j h�@������p���j �E�P�����Q�M��"�������������������������������t�M�e����M������E�9j�E�P�M��դ��j�j��EP�M�Q�M��ͬ���E�P�M�h����M�跚���ER��P�h�#���XZ_^[��,  ;��l�����]Ë�   p����   �����   �str pos ����������������������������������������������������������������������������������������������������������������U���P  SVW�������T   ������EP�PX螗��P�M��i���j h�@����������j �E�P������Q�M�薰�������������������聙����������t�M�ٰ���M��f����E�>  j�E�P�M��F���j�j��EP�M�Q�M��>���j h�@�������`���j �E�P������Q�M�����������������������������������t�M�U����M������E�   j�E�P�M��¢��j�j��EP�M�Q�M�躪��j h�@������ܲ��j �E�P�����Q�M�莯�������������������y�����������t�M�ѯ���M��^����E�9j�E�P�M��A���j�j��EP�M�Q�M��9����E�P�M�Բ���M��#����ER��P��菜��XZ_^[��P  ;��ت����]Ë�   ����    ����   str pos ��������������������������������������������������������������������������������������������������������������������������������������������U���t  SVW�������]   ������EP�PX����P�M�蹱��j h�@�������4���j �E�P������Q�M�����������������������і����������t�M�)����M�趖���E��  j�E�P�M�薠��j�j��EP�M�Q�M�莨��j h�@������谰��j �E�P������Q�M��b���������������������M�����������t�M襭���M��2����E�>  j�E�P�M�����j�j��EP�M�Q�M��
���j h�@�������,���j �E�P������Q�M��ެ��������������������ɕ����������t�M�!����M�讕���E�   j�E�P�M�莟��j�j��EP�M�Q�M�膧��j h�@�����訯��j �E�P�����Q�M��Z��������������������E�����������t�M蝬���M��*����E�9j�E�P�M�����j�j��EP�M�Q�M������E�P�M蠯���M������ER��P�0�[���XZ_^[��t  ;�褧����]Ë�   8����   T����   Pstr pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������EP�DX�Q<�B�Ѓ�;�肦��_^[���   ;��r�����]���������������������������������U���p  SVW�������\   ������ǅ����    j h�>�������q���P�ɕ�����E��������$����}� u3���   �E�    �E�P�M�� ����E�P�M�Q�M����������   �}���   �M��o����E��}� tF�EP�������-���������Pj������Q�M��6�����������訔����tǅ����   �
ǅ����    ��������������������t��������������X�����������t��������������;�����������t�EԉE�������E�R��P��菖��XZ_^[��p  ;��ؤ����]Ë�   ����   3����   /����   (browse dat id ��������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�訐�������_^[���   ;��أ����]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bx��;��}���_^[���   ;��m�����]� �������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R�DX�P�M����   ��;�� ���P�M�Ǫ���� ��������E_^[���   ;��٢����]� �������������������������������������U���d  SVW�������Y   ������ǅ����    �} u6j h�>�������˩��P�#������E�������~����} u3��$  �E�    �EP�M��z����E�P�M�Q�M��O�������   �}���   �M��ɕ���Eă}� tF�EP������臦��������Pj������Q�M�萧����������������tǅ����   �
ǅ����    ��������������������t�������������貎����������t�������������蕎����������t�E��E��2�+�}�u%�}� t�EP�M��5������n�����t�E��E��������E�R��P��輒��XZ_^[��d  ;�������]ÍI    �����   ����   ����   �browse dat id ��������������������������������������������������������������������������������������������������������������������������������������U����   SVW������:   ������} u3��   �EP�M��J����E�    �E�    �E�P�M�Q�M�������tT�}�t�}�u"�EP�M�艓��P�ה������t�   �*�$�}�u�EP�M�虍�����Ҏ����t�   ��3�R��P�d�%���XZ_^[���   ;��n�����]�   l����   �����   �����   �dat id browse ����������������������������������������������������������������������������������U����   SVW��@����0   ������DX�H<��Q��;�語��_^[���   ;�蚞����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �@�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M�轓���E��t�E�P�ɏ�����E�_^[���   ;��ܝ����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �@_^[��]��������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;�����������
ǅ���    �E�    _^[���   ;�������]������������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M���  ��;�����_^[���   ;��o�����]������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M���(  ��;�����_^[���   ;��������]������������������������������U����   SVWQ������<   ������Y�M������P�DX�Q�M���   ��;�藛��P�M讣��������h����E_^[���   ;��p�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M���$  ��;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�DX�B��  �у�;�苚��_^[���   ;��{�����]��������������������������U����   SVW��@����0   �������EP�DX�Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   ������DX�H��  ��;�跙��_^[���   ;�觙����]����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��H���_^[���   ;��8�����]�����������������������U����   SVW��@����0   �������EP�MQ�DX�B��x  �у�;��ۘ��_^[���   ;��˘����]��������������������������U����   SVW��@����0   �������EP�DX�Q��|  �Ѓ�;��o���_^[���   ;��_�����]������������������������������U����   SVW��@����0   ������DX�H��d  ��;�����_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ�DX�B��p  �у�;�蛗��_^[���   ;�苗����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B��t  �у�;��+���_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M��M��e�����E�P�DX�Q$�BD�Ѓ�;�赖���E�_^[���   ;�袖����]���������������������������������U����   SVWQ��4����3   ������Y�M��M�������E�P�DX�Q$�BD�Ѓ�;��5�����EP�M�Q�DX�B$�Hd�у�;������E�_^[���   ;�� �����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��5�����E�P�DX�Q$�BD�Ѓ�;�腕����EP�M�Q�DX�B$�H�у�;��c����E�_^[���   ;��P�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M�腙����E�P�DX�Q$�BD�Ѓ�;��Ք����E�P�MQ�DX�B$�HL�у�;�賔���E�_^[���   ;�蠔����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q$�BH�Ѓ�;��-����M��L���_^[���   ;�������]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�HL�у�;�詓��_^[���   ;�虓����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q$�M��B��;��!���_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q$�M��Bl��;�譒��_^[���   ;�蝒����]� �������������������������U����   SVWQ��4����3   ������Y�M��DX�P$��M��Bp��;��B���_^[���   ;��2�����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q$�B�Ѓ�;��͑��_^[���   ;�轑����]����������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q�DX�B$�H�у�;��V���P�M������ ����i~���E_^[���   ;��/�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H�у�;�蹐��_^[���   ;�詐����]� �������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q�DX�B$�H �у�;��6���P�M�M�������������E_^[���   ;�������]� �������������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q�DX�B$�H$�у�;�薏��P�M譗��������g����E_^[���   ;��o�����]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M���������{��������ہ���E_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q$�B(�Ѓ�;��}���_^[���   ;��m�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�DX�Q$�Bh�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H,�у�;�虍��_^[���   ;�艍����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H0�у�;�����_^[���   ;��	�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H4�у�;�虌��_^[���   ;�艌����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H8�у�;�����_^[���   ;��	�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�DX�B$�HL�у�;�虋���E�_^[���   ;�膋����]� ����������������������������������U����   SVW������9   ������EP�M��T�����EP�M�Q�DX�B$�H@�у�;������E�P�M�&����M���}���ER��P��-�|��XZ_^[���   ;��ڊ����]�    .����   .fn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H@�у�;��I����E�_^[���   ;��6�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H<�у�;��ɉ��_^[���   ;�蹉����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�H<�у�;��I��������_^[���   ;��2�����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H$�QP�҃�;��ƈ��_^[���   ;�趈����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B$�HT�у�;��I���_^[���   ;��9�����]� �������������������������������������U����   SVW��@����0   ������DX�H$��QX��;��ڇ��_^[���   ;��ʇ����]�������������������������U����   SVW��@����0   �������EP�DX�Q$�B\�Ѓ�;��r���_^[���   ;��b�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q$�B`�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVW��@����0   ������DX�H(����;�苆��_^[���   ;��{�����]��������������������������U����   SVW��@����0   �������E�Q�DX�B(�H�у�;�� ����E�     _^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�DX�P(�M��B��;�芅��_^[���   ;��z�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P(��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��B��;�蝄��_^[���   ;�荄����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P(�M��B��;��&���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B(�M��P ��;�詃��_^[���   ;�虃����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ�DX�B(�M��P��;��'���_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P(�M��B$��;�覂��_^[���   ;�薂����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��DX�P(��M��B(��;��2���_^[���   ;��"�����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P(��M��B,��;����_^[���   ;�貁����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P(��M��B0��;��R���_^[���   ;��B�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��B4��;��݀��_^[���   ;��̀����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��BX��;��m���_^[���   ;��]�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��B\��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��B`��;����_^[���   ;��}����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bd��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bh��;��~��_^[���   ;��~����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bl��;��=~��_^[���   ;��-~����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bx��;���}��_^[���   ;��}����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M����   ��;��Z}��_^[���   ;��J}����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bt��;���|��_^[���   ;���|����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��Bp��;��}|��_^[���   ;��m|����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��r����t2�M��Q�M��r����t�U��R�M���q����tǅ0���   �
ǅ0���    ��0���_^[���   ;���{����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��p�����t8�MQ�A�$�M��Z�����t"�UQ�B�$�M��D�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��{����]� ������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��2z����t2�M��Q�M��z����t�U��R�M��z����tǅ0���   �
ǅ0���    ��0���_^[���   ;��Yz����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M���m����t<�M���A�$�M���m����t$�U���B�$�M��m����tǅ0���   �
ǅ0���    ��0���_^[���   ;��y����]� ����������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M���t����tE�M��Q�M���t����t2�U��R�M��t����t�E��$P�M��t����tǅ0���   �
ǅ0���    ��0���_^[���   ;���x����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��r����tE�M��Q�M��pr����t2�U��R�M��]r����t�E��$P�M��Jr����tǅ0���   �
ǅ0���    ��0���_^[���   ;���w����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��`����tE�M��Q�M��`����t2�U��0R�M��`����t�E��HP�M��r`����tǅ0���   �
ǅ0���    ��0���_^[���   ;��&w����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��L�����tE�M��Q�M��9�����t2�U��0R�M��&�����t�E��HP�M�������tǅ0���   �
ǅ0���    ��0���_^[���   ;��Vv����]� ��������������������������������������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M���`����u3���   �}� u)������Wz��P�M�f���������b���   �   ��h�@��@��P�M�Q�DX�B���   �у�;��xu���E��}� uj��M��(v��3��Lj �E�P�M�Q�M��]b����u�E�P�n����3��&j �E��P�M�Q�M�v���E�P�~n�����   R��P��C�f��XZ_^[���   ;���t����]�    �C����   D����    Dc len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�DX�Q�B�Ѓ�;��!t��_^[���   ;��t����]� �����������������������������U����   SVWQ������?   ������Y�M��M��Ux���E�P�M��m����uǅ���    �M���`��������$�E�P�M�A`��ǅ���   �M��`�������R��P��E�e��XZ_^[���   ;��Ts����]�    �E����   �Estr ��������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�P�M��g����u3���E�����؋M��   R��P�DF�Id��XZ_^[���   ;��r����]� ��   LF����   XFc ��������������������������������������U����   SVWQ��4����3   ������Y�M��} ����Q�M��#{��_^[���   ;��r����]� ��������������������U����   SVWQ������=   ������Y�M�j �M�j�����E���h�@��@��P�M�Q�DX�B���   �у�;��q���Eԃ}� uj��M��<r��3��dj �E�P�M�Q�M�u���E�P�M��m`����t �M�Q�U�R�M���w����tǅ���   �
ǅ���    ������E�E�P�xj�����E�R��P��G�b��XZ_^[���   ;���p����]�    �G����   �Gmem ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bd��;��=p��_^[���   ;��-p����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�DX�P�M��Bh��;���o��_^[���   ;��o����]� ����������������������������������U����   SVWQ������<   ������Y�M��� ���P�M�L\��P�M��by��������� ����i\�������_^[���   ;��,o����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q(�M��B8��;��n��_^[���   ;��n����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q(�M��B<��;��Ln��_^[���   ;��<n����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q(�M��B@��;���m��_^[���   ;���m����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q(�M��BD��;��lm��_^[���   ;��\m����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��BH��;���l��_^[���   ;���l����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B(�M��P|��;��l��_^[���   ;��yl����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q(�M��BL��;��l��_^[���   ;���k����]� �������������������������U����   SVWQ��4����3   ������Y�M�����E�$�DX�P(�M��BT��;��k��_^[���   ;��k����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�DX�P(�M��BP��;��k��_^[���   ;��k����]� �����������������������U����   SVW��@����0   ������DX�H(��Q��;��j��_^[���   ;��j����]�������������������������U����   SVW��@����0   �������E�Q�DX�B(�H�у�;��Pj���E�     _^[���   ;��7j����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�DX�Q(�M����   ��;��i��_^[���   ;��i����]�( ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�DX�B(�H�у�;��"i��_^[���   ;��i����]���������������������������������U����   SVW��@����0   ������DX�H,��Q,��;��h��_^[���   ;��h����]�������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B4��;��Rh��_^[���   ;��Bh����]���������������������������������U����   SVW��@����0   �������E�Q�DX�B,�H0�у�;���g���E�     _^[���   ;���g����]��������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B8��;��bg��_^[���   ;��Rg����]���������������������������������U����   SVWQ������<   ������Y�M������P�DX�Q,�M��B<��;���f��P�M�o��������Y���E_^[���   ;���f����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q�DX�B,�M��P@��;��Vf��P�M�n���� ����iS���E_^[���   ;��/f����]� �������������������������������������������U����   SVW��@����0   �������j j �DX�H,��҃�;���e��_^[���   ;��e����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H,�Q�҃�;��Fe��_^[���   ;��6e����]� ����������������������������������U����   SVW��@����0   �������E�Q�DX�B,�H�у�;���d���E�     _^[���   ;��d����]��������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B��;��Rd��_^[���   ;��Bd����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B��;���c��_^[���   ;���c����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B��;��rc��_^[���   ;��bc����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B ��;��c��_^[���   ;���b����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B$��;��b��_^[���   ;��b����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P,��M��B(��;��"b��_^[���   ;��b����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B,�M��P��;��a��_^[���   ;��a����]� �������������������������������������U����   SVWQ������<   ������Y�M������P�DX�Q,�M��B��;��*a��P�M�Ai���������S���E_^[���   ;��a����]� �������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��D  �҃�;��`��_^[���   ;��`����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��H  �҃�;��(`��_^[���   ;��`����]�����������������������U����   SVW��@����0   �������EP�DX�Q��L  �Ѓ�;��_��_^[���   ;��_����]������������������������������U����   SVW��@����0   �������EP�MQ�DX�B�H�у�;��N_��_^[���   ;��>_����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H�Q�҃�;���^��_^[���   ;���^����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B�H�у�;��n^��_^[���   ;��^^����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H�Q�҃�;���]��_^[���   ;���]����]��������������������������U����   SVW��@����0   �������EP�MQ�DX�B�H�у�;��]��_^[���   ;��~]����]�����������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;��]��_^[���   ;��]����]��������������������������U����   SVW��@����0   �������EP�DX�Q�B�Ѓ�;��\��_^[���   ;��\����]���������������������������������U���  SVW�������E   ������E�P�M�IN���M��E����uǅ����    �M��O���������   j�E�P�S������u*�E�P�f`������uǅ����    �M���N���������Tj�EP��R������u*�EP�:_������uǅ���    �M��N��������ǅ���   �M��N�������R��P�X]�1M��XZ_^[��  ;��z[����]�   `]����   l]parent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP�DX�Q�B �Ѓ�;���Z��_^[���   ;���Z����]���������������������������������U����   SVW��@����0   �������EP�MQ�DX�B�H(�у�;��^Z��_^[���   ;��NZ����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�DX�B��  �у�;���Y��_^[���   ;���Y����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q��   �Ѓ�;��cY��_^[���   ;��SY����]����������������������������������U����   SVW��@����0   �������EP�DX�Q��  �Ѓ�;���X��_^[���   ;���X����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H��  �҃�;��xX��_^[���   ;��hX����]�����������������������U����   SVW������9   ������� ���P�DX�Q�B$�Ѓ�;��X��P�M�&`���� �����J���E_^[���   ;���W����]���������������������������������������U����   SVW������9   ������� ���P�DX�Q���  �Ѓ�;��|W��P�M�_���� ����MJ���E_^[���   ;��UW����]������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;���V��_^[���   ;���V����]��������������������������U���$  SVW�������I   ������ǅ8���    �=,] t!������P�,]�pH����8����������������\����8���������������������������R�M�Y^����8�����t��8����������I����8�����t��8������������H���E_^[��$  ;���U����]�����������������������������������������������������������U����   SVW������9   �������EP�� ���Q�DX�B���  �у�;��hU��P�M�]���� ����9H���E_^[���   ;��AU����]��������������������������������U����   SVW��@����0   ������j�EP��X�����E_^[���   ;���T����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��xT��_^[���   ;��hT����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��T��_^[���   ;���S����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��S��_^[���   ;��S����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�DX�H���  �҃�;��(S��_^[���   ;��S����]�����������������������U����   SVW��@����0   ������DX�H���   ��;���R��_^[���   ;��R����]����������������������U����   SVW��@����0   �������EP�DX�Q���   �Ѓ�;��_R���E�     _^[���   ;��FR����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M����;���Q��_^[���   ;���Q����]� ������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M��B��;��bQ��_^[���   ;��RQ����]���������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;���P��_^[���   ;���P����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B`��;��}P��_^[���   ;��mP����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bd��;��P��_^[���   ;���O����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bh��;��O��_^[���   ;��O����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bl��;��-O��_^[���   ;��O����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bp��;��N��_^[���   ;��N����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bt��;��MN��_^[���   ;��=N����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���M��_^[���   ;���M����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M���  ��;��jM��_^[���   ;��ZM����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��Bx��;���L��_^[���   ;���L����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��L��_^[���   ;��zL����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B|��;��L��_^[���   ;��L����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��K��_^[���   ;��K����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��:K��_^[���   ;��*K����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���J��_^[���   ;��J����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��ZJ��_^[���   ;��JJ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���I��_^[���   ;���I����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��zI��_^[���   ;��jI����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��
I��_^[���   ;���H����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��H��_^[���   ;��H����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��*H��_^[���   ;��H����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��G��_^[���   ;��G����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��  �у�;��FG��_^[���   ;��6G����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;���F��_^[���   ;��F����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;��FF��_^[���   ;��6F����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���E��_^[���   ;��E����]� ����������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q�DX�B �H$�у�;��SE����tǅ0���   �
ǅ0���    ��0���_^[���   ;��#E����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR�DX�H �QL�҃�;��D��_^[���   ;��D����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q�DX�B �H(�у�;��D���   _^[���   ;��
D����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q�M��B��;��C��_^[���   ;��C����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q�M��B��;��,C��_^[���   ;��C����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q�M��B��;��B��_^[���   ;��B����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�DX�Q�M��B��;��LB��_^[���   ;��<B����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B��;���A��_^[���   ;���A����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B��;��mA��_^[���   ;��]A����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M��P\��;���@��_^[���   ;���@����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M���  ��;��v@��_^[���   ;��f@����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�DX�P�M��B ��;���?��_^[���   ;���?����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�DX�P�M��B$��;��{?��_^[���   ;��k?����]� �����������������������U����   SVWQ��4����3   ������Y�M�����E�$�DX�P�M��B(��;��	?��_^[���   ;���>����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B,��;��>��_^[���   ;��}>����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B0��;��>��_^[���   ;��>����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B4��;��=��_^[���   ;��=����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B8��;��==��_^[���   ;��-=����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B<��;���<��_^[���   ;��<����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��B@��;��]<��_^[���   ;��M<����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��BD��;���;��_^[���   ;���;����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��BH��;��};��_^[���   ;��m;����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��BL��;��;��_^[���   ;���:����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��BP��;��:��_^[���   ;��:����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M����   ��;��:��_^[���   ;��:����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M��BT��;��9��_^[���   ;��9����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�DX�B��  �у�;��69��_^[���   ;��&9����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M����   ��;��8��_^[���   ;��8����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�DX�Q�M����   ��;��.8��_^[���   ;��8����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M��PX��;��7��_^[���   ;��7����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;��?7��_^[���   ;��/7����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���6��_^[���   ;��6����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;��Z6��_^[���   ;��J6����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�DX�Q�M����   ��;���5��_^[���   ;���5����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;��v5��_^[���   ;��f5����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;���4��_^[���   ;���4����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�DX�B�M����   ��;��4��_^[���   ;��v4����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;��4��_^[���   ;���3����]������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;��3��_^[���   ;��3����]������������������������������U����   SVWQ��4����3   ������Y�M��DX�P��M����   ��;��/3��_^[���   ;��3����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�DX�B���   �у�;��2��_^[���   ;��2����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�DX�Q��   �Ѓ�;��32��_^[���   ;��#2����]����������������������������������U����   SVW��(����6   �������EP�MQ��,���R�DX�H���  �҃�;��1��P�M�|9����,��������E_^[���   ;��1����]���������������������������������������������U����   SVW��@����0   �������EP�MQ�DX�B���  �у�;��1��_^[���   ;��1����]��������������������������U����   SVW��4����3   ������j�   ���E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;��0��_^[���   ;��o0����]����������������������������������������������U����   SVW��@����0   ������hdX�EPh�f �E����_^[���   ;���/����]�������������������������U����   SVW������<   ������j�{������E��}� t	�E��x uǅ��������M�w"��������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�7���EP�M��Q�҃�4�� ����M�0"���� ���_^[���   ;��5/����]����������������������������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;��.��_^[���   ;��.����]�����������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�M��Q�҃�;��.��_^[���   ;��.����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� (A�M��N��_^[���   ;��-����]�������������������������U����   SVWQ��4����3   ������Y�M��M��D(���E��t�E�P������E�_^[���   ;��,-����]� ������������������������U����   SVWQ��(����6   ������Y�M��M����E�M��Q�P�E�M��Q�P�E�    �	�E���E�E��M�;H}�E��H�U��P�M� ����u3���͸   _^[���   ;��z,����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��} |$�E��M;H}�} |�E��M;H}�E;Eu�"�E��H�U��P�M��Q�E��Q������_^[���   ;���+����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E;E}	�E���E�} |$�E��M;H}�} |�E��M;H}�E;Eu�/�E��H�U���E�EP�M������t�EP�M�Q�M����_^[���   ;���*����]� �������������������������������������������U����   SVWQ������9   ������Y�M��E��x u�E��H�M��%�E��x t�E��H�U�J�M���E��H��M��}� u3��]��h0A��@��P�M���Q�U��BP�DX�Q��  �Ѓ�;��/*���E�}� u3���E��M�H�E��M��H�   _^[���   ;���)����]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��P;Qu�M���"����u3��&�E��H�U��B�U���E��H���U��J�   _^[���   ;��G)����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��M;H}�EP�MQ�M��j&���#�E��H;M}j �M�������EP�M����_^[���   ;��(����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3���E��H�U�E���   _^[��]� ���������������������������U����   SVWQ��(����6   ������Y�M��E��M;H~	�E��H�M�} }�E    �E��M��P;Qu�M��)!����u3��Z�E��H�M��	�E���E�E�;E~�E��H�U��B�U�u�L�����ԋE��H�U�E���E��H���U��J�   _^[���   ;��B'����]� ��������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3��E�E��H���U��J�	�E���E�E��M;H}�E��H�U��B�U�u�L����Ѹ   _^[��]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����P�M����_^[���   ;��&����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E��M�;H}�E��H�U��;Eu�E���ԃ��_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��E���P������E��@    �E��@    �M��A    _^[���   ;���$����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��@    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M��E��H��Q�M�����E�}� t�E��H��Q�M��.���E�_^[���   ;��+$����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H}�E��H�U���3�_^[��]� �������������������U����   SVWQ��$����7   ������Y�M��EP�M��T��j�E��HQ�U��BP�M��~��R��P�������XZ_^[���   ;��F#����]� ��   ������   ��sort ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��*���E�� �A�E��M�H�E�_^[���   ;��"����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�Ѓ�;��O"��_^[���   ;��?"����]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�� �A�E�_^[��]���������������������������U����   SVWQ��$����7   ������Y�M��EP�M��t��j�E��HQ�U��BP�MQ�M��)��R��P�t����XZ_^[���   ;��b!����]� ��   |�����   ��sort �����������������������������������U����   SVWQ��4����3   ������Y�M��E�� �A�M�����'���M�����'���E��@    �M�����E�_^[���   ;�� ����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �A�E��@    �E��@    �E�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��M��!*���E��t�E�P�������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�����E��t�E�P�Y�����E�_^[���   ;��l����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� �A�M��$���M����-)���M����")��_^[���   ;�������]�����������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E����M��A�E����M��A�E��@    _^[��]���������������������������U���   SVWQ�� ����@   ������Y�M��M���$���E��}� tm�M��v)���E�}� tM�E��������������������� t%��j��������������;������� ����
ǅ ���    �E�    �E�E�덋M����_^[��   ;������]����������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t�M��Q�z t�E��H��0����
ǅ0���    ��0���_^[��]������������������������������������U����   SVWQ��0����4   ������Y�M��E����M�9At�U��B��0����
ǅ0���    ��0���_^[��]���������������������������U����   SVWQ������9   ������Y�M��M��#���E��}� t�M��'���E�M��U!���E�E���_^[���   ;������]������������������������������U����   SVWQ������:   ������Y�M��E�    �M��"���E��}� tD�E�M�U���U�;�uǅ���   �
ǅ���    ����� t�E���M���&���E��3�_^[���   ;��m����]� �����������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E�M��Q�P�E����M�A�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E����M�A�E�M��Q�P�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ������9   ������Y�M��E�    �M��� ���E���M��S%���E��}� t�E���E���E�_^[���   ;�������]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �A�M����_^[���   ;��j����]�������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t;�E��x t2�E��H�U��B�A�E��H�U��B�A�E��@    �M��A    _^[��]�����������������������������������U����   SVW��4����3   ������E��M��E�M���E�M��_^[��]������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ�����_^[���   ;������]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�`	�����E��}� u3��5�M��
���E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;��+����]������������������������������������������U����   SVWQ������9   ������Y�M���EP�DX�Q�M��Bd��;�����E�}� u3��s��h�A�PA��P�M��Q�DX�B���   �у�;��~���E��}� u3��4��EP�M��Q�U�R�DX�P�M��Bh��;��I���E�E��  �E�_^[���   ;��-����]� ���������������������������������������������������������U����   SVW��@����0   ������j h�  hhX�M�h���hX_^[���   ;������]����������������������U����   SVW��@����0   ������j h�  hhX�M����hX_^[���   ;��G����]����������������������U����   SVW��@����0   ������h� �M�E	����tj h�  hhX�M�A	��������hBhhX�������hX_^[���   ;������]������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�DX���   �M��B��;��J��_^[���   ;��:����]� ����������������������U����   SVWQ��4����3   ������Y�M��DX���   ��M��Bx��;�����_^[���   ;�������]������������������������������U����   SVW��(����6   ������j h�  hhX��,���P�M�e����������,��������hX_^[���   ;��N����]�����������������������������U����   SVW��(����6   ������j h�  hhX��,���P�M������������,����
����hX_^[���   ;�������]�����������������������������U���  SVW�������B   �����󫡐A3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |I�E�M������E��E���
}�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�먋E��D� j �E�P�M�=���ER��P� ��s��XZ_^[�M�3��������  ;������]�   (�����   4�hexstring ����������������������������������������������������������������������������������U���  SVW��x����b   ������} ��   �}   @��   j h4B�������R��Pj0j jj �E�U��������x�����|���߭x����5(B���$������P�������P�MQ�Z���������������������������E�^  �  �} ��   �}   ��   j h B���������Pj0j jj �E�U�
�R�����x�����|���߭x����5(B���$������P�T�����P�MQ�������������#��������������E��   �r�} |l	�}   vaj hB�������!��Pj0j jj �m�5(B���$������P�������P�MQ�E��������������������������E�Lj hB���������P�EP��,���Q�.����P�UR���������,����^���������S����E_^[�Ĉ  ;������]��������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��(����6   �������EP��,���Q�DX�B�H(�у�;��;��P�M�����,����N����E_^[���   ;������]�����������������������������������U����   SVW��(����6   ��������E P�MQ�UR�EP���E�$��,���Q�DX�B�H$�у�;����P�M�\����,��������E_^[���   ;��n����]���������������������������������������������U����   SVWQ��0����4   ������Y�M��E�M��;t3���   �E�x uN�E�8 uF�E�x u=�E��x u�M��9 u�U��z uǅ0���   �
ǅ0���    ��0����   �R�E��x uI�E��8 uA�E��x u8�E�x u�M�9 u�U�z uǅ0���   �
ǅ0���    ��0����M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� �������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����������_^[���   ;��h
����]� ��������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M���	���8 t��E�_^[���   ;���	����]����������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M��L	���8 t(�E�P�M�;	��P�M�Q�M��.	�����D����t�뾃} t�E�M��}� ~�E�P�M������8 uǅ$���   �
ǅ$���    ��$���_^[���   ;��	����]� �����������������������������������������������������������U����   SVW��4����3   ������j�k   ���E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;��p��_^[���   ;��`����]�������������������������������U����   SVW��@����0   ������h]�EPhD �E�����_^[���   ;�������]�������������������������U����   SVWQ��(����6   ������Y�M�j\�v������E�}� t	�E�x\ u���E�P�M�Q\�҃�;�����E�_^[���   ;��r����]���������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;������EP�M�������E�_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�F������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��U���EP�M��n����E�_^[���   ;��6����]� ����������������������������������U����   SVWQ������;   ������Y�M�j\�������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;�����EP���������P�M�������E�_^[���   ;������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U����   SVWQ��(����6   ������Y�M�j\�������E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;�����EP�M������EP�M�������E�_^[���   ;��z����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;������EP�M������EP�M��#����EP�M������E�_^[���   ;������]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�&������E�}� t	�E�x` u���E�P�M�Q`�҃�;��5��_^[���   ;��%����]������������������������������������U����   SVWQ��(����6   ������Y�M�jd�������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jl�v������E�}� t	�E�xl u���E�P�M�Ql�҃�;����_^[���   ;��u����]������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��� ��_^[���   ;��� ����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��F ��_^[���   ;��6 ����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u�]���EP�M�Q�U�Bp�Ѓ�;�����_^[���   ;�������]� ����������������������������������������U����   SVWQ������:   ������Y�M�jt�������E�}� t	�E�xt uh]�M�|����E�:��EP�M�Q�����R�E�Ht�у�;������P�M��������������E_^[���   ;��������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�jx�6������E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;��>����E�_^[���   ;��+�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j|�������E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j|��������E�}� t	�E�x| u�   �#��E�P�MQ�U�B|�Ѓ�;�����������_^[���   ;��������]� ���������������������������������U����   SVWQ������:   ������Y�M�h�   �S������E�}� t�E샸�    u�E��4��EP�M�Q�����R�E싈�   �у�;��N�������������E�_^[���   ;��0�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��4����3   ������j�[������E��}� t	�E��x u3���E���H��;��o���_^[���   ;��_�����]������������������������������U����   SVW��4����3   ������E�8 u�?j��������E��}� t	�E��x u�!��EP�M��Q�҃�;�������E�     _^[���   ;��������]��������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j�,������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;��1���_^[���   ;��!�����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;�����_^[���   ;�������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;������_^[���   ;��������]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j �F������E�}� t	�E�x  u3����E�P�M�Q �҃�;��S���_^[���   ;��C�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j$�������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;������_^[���   ;�������]����������������������������������U����   SVWQ��(����6   ������Y�M�j(�&������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;��'���_^[���   ;�������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;�����_^[���   ;��{�����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;������_^[���   ;��������]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j4�F������E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��S���_^[���   ;��C�����]����������������������������������U����   SVWQ��(����6   ������Y�M�j8�������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;�����_^[���   ;�������]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�������E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��(����6   ������Y�M�jD�v������E�}� t	�E�xD u3����E�P�M�QD�҃�;�����_^[���   ;��s�����]����������������������������������U����   SVWQ��(����6   ������Y�M�jH��������E�}� u���EP�M�Q�U�BH�Ѓ�;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jL�V������E�}� u3����EP�M�Q�U�BL�Ѓ�;��h���_^[���   ;��X�����]� ������������������������������������U����   SVWQ��(����6   ������Y�M�jP��������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;������_^[���   ;��������]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�6������E�}� u3����E�P�M�QT�҃�;��L���_^[���   ;��<�����]���������������������������U����   SVWQ��(����6   ������Y�M�jX�������E�}� u���EP�M�Q�U�BX�Ѓ�;������_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;��"���_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��z���_^[���   ;��j�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;������_^[���   ;��������]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �C������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��R���_^[���   ;��B�����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;������_^[���   ;�������]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��,���_^[���   ;�������]� ����������������������������������������U����   SVW������9   ������h�   �������E��}� u�M�D����E�9��EP�� ���Q�U����   �Ѓ�;�����P�M�R����� ��������E_^[���   ;��d�����]���������������������������������������������������U����   SVW��$����7   ������h�   ��������E��}� t�E����    u�EP�M�}����E�=��EP�MQ��(���R�E����   �у�;�����P�M�I�����(����x����E_^[���   ;�������]�����������������������������������������������U����   SVWQ������?   ������Y�M�h�   ��������E�}� t�E샸�    uj ����������P�M�]����E�9��EP�����Q�U�M����   ��;������P�M�n�������������E_^[���   ;�������]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;�����_^[���   ;�������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�U�M����   ��;��j���_^[���   ;��Z�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�U�M����   ��;������_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����EP�U�M����   ��;��*���_^[���   ;�������]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����E�M����   ��;�����_^[���   ;��~�����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;������_^[���   ;��������]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u���EP�U�M����   ��;��<���_^[���   ;��,�����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;�����_^[���   ;�������]� ����������������������������������������������U����   SVWQ������9   ������Y�M�h�   ��������E�}� t�E샸�    u3����E�M����   ��;�������E��E�_^[���   ;��������]���������������������������������������U����   SVWQ��(����6   ������Y�M���E�P�DX���   �BX�Ѓ�;��j����E�}� u3���EP�MQ�M��h���_^[���   ;��=�����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H|�Q�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P�DX���   �BX�Ѓ�;��J����E�}� u3���EP�MQ�M��@���_^[���   ;�������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�DX�H|�Q8�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q�DX�B�H�у�;������U��B�E�_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q�DX�B�H�у�;������U��B_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��E��HQ�UR�EP�M��R�DX�H�Q�҃�;�� ����M��A�   _^[���   ;��������]� ���������������������������������U����   SVW��<����1   ������E��<�����<���t��E�4]�E�0]�   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$�L��   �]  �8]���8]�=8]��   �EP������=�2  }
������&  �} u
������  h8B�TA��Ph?]j��������� ����� ��� t�� �������������
ǅ���    ������,]�=,] t�EP�,]�j����   �   �EP�MQ���������u����   �   �|�	����u�8]���8]u\�����,����=,] t?�,]��8�����8�����,�����,��� tj��,�������������
ǅ���    �,]    �   ����_^[���   ;�������]Ð��������4�������������������������������������������������������������������������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�������}�EP�M�Q�U�R�M���������U��������_^[��,  ;��n�����]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M�������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��<�����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�������}�E�P�M�Q�U�R�M���������U��������_^[��8  ;��������]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M�������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;�������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��[�����}�E�P�M�Q�U�R�M��
������U��������_^[��8  ;��%�����]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��u�EP�MQ�UR�M��v����83��} ����t�EP�MQ�UR�M��������EP�MQ�UR�M��Q���_^[���   ;�������]� �������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  �Ek� E�E���E�P�MQ�U���M����;�������Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;��r����Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��0�����t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;��������]� ����������������������������������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u�E� ����3���  �Ek� E�E���E�P�MQ�U���M����;��
����Eȃ}� u
�E��  ��}� }�E�     3��  �E�   �E���E��E�    �E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;������Eȃ}� uS�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��G�����t�
��E��E�뷋E���   ��}� }�Eԃ��E��	�Eԃ��E��D����}� ~�Eԃ��M���E�Mԉ�E�;M}F�E�M�M�M���E�P�MQ�U���M����;�������|h�B�XA��9P�|������E�8 ~I�E����MM�M���E�P�MQ�U���M����;��l�����h�B�XA��?P�+�����3�_^[��  ;��@�����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������u�U��� PRSVW�Ej P�;�����_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR�b������E�@���E�;|�_^[��]���������������������������̋�U��V���t!��tS�]��tW�̋�����F�V�3_[^]� �������������̋�U��QSVW��3���;�tR�}�9>~K��    �F�8�����9T�u�D8�9t�N�T�ERP����������̋E�@���E�;|������̋u3��ƅ�tV�@G��u���tJ9u9Vu
9Vu9Vt�MWVQ�8���������̋F9T0�t�MWVQ����������̋vO��u�_^[��]� �����������������������������������������������������������̀=@] uj jj j j �@]�����P������������������������������jjj j j ��������������������̋�U���4����} t舵����]�������̋�U����A����AO���A���A���A���A����Ag���A����A����A�]�������������������������������������̋�U��Q�D]�E��M�D]�E���]������������������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������������������������������������������������������̋�U��Q�M��EP�M�Q���������]� ����������������̋�U��Q�M��E�� �B�M�Q课������]��������������̋�U��Q�M��M��8����E��t�M�Q�ӽ�����E���]� �����������������̋�U��Q�M��EP�M�Q��������]� ����������������̋�U��Q�M��E�P�e�������]�������̋�U��Q�M��E���	P�M��	Q�8������������]� �������������������̋�U��Q�M��E���	P�M��	Q�����������؋�]� ��������������������̋�U��Q�M��E���	P�M��	Q踾����3҅���]� �����������������̋�U��Q�M��E�����]�������������̋�U��Q�M��E�� �B�E���]� ��������������������̋�U��Q�M��E���]� �������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������������̋�U��j�h`+h�d�    P���SVW��A1E�3�P�E�d�    �}��   �`�����u3��  �������u����3��  ����������������L]�H�����}�?���讽��3��i  �J�����|�������|j �o�������t�����	����x���3��3  j�S������H]���H]�  �} um�=H] ~X�H]���H]�E�    �=�] u�^����������������E������   ��} u�=�A�t�}�����3��   �   �}��   �����h�   h�Bjh  j�)������E�}� tV�U�R��AP��]Q�ܑ�Ѕ�t%j �U�R��������ؑ�M��U��B�����j�E�P�f�����3���3����}u
j �y������   �M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��}u�P����EP�MQ�UR�   ��]� �����������������������̋�U��j�h�+h�d�    P���SVW��A1E�3�P�E�d�    �e��E�   �} u�=H] u3��N  �E�    �}t�}uT�=�B t�EP�MQ�UR��B�E�}� t�EP�MQ�UR�l����E�}� u�E�    �E������E���   �EP�MQ�UR������E�}u=�}� u7�EPj �MQ�۲���URj �EP�����=�B t�MQj �UR��B�} t�}u@�EP�MQ�UR�������u�E�    �}� t�=�B t�EP�MQ�UR��B�E��E������8�E���U��E�P�M�Q�׽����Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������̋T$�L$��ti3��D$��u���   r�=�� t�X���W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̋�U��Qj j j�@_P�MQ�R������E��E���]������������������������̋�U��j�EP�P�����]������������;�Au����������������������̋�U��j�h�+h�d�    P���SVW��A1E�3�P�E�d�    �`����E�    �EP�Y   ���E��E������   ��N���ËE�M�d�    Y_^[��]������������������������������������������̋�U������P�ܑ�E����Q�ܑ�E��U�;U�r�E�+E�����s3���   j�M�Q��������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}h8Cj�E�P�M�Q��������E��}� u:�U���U�E�;E�r%h�   h8Cj�M�Q�U�R�������E��}� u3��Q�E�+E����M����U��E��E��M�Q������UR���M���U����U��E�P������E��]�����������������������������������������������������������������������������������������������̋�U��EP����������؃�]��������������������̋�U��Qh�   h8Cjjj ��������E��E�P������������}� u�   ��U��    3���]������������������������̋�U��Q�tjP�ܑ�E��}� t�U�j�������jj �֭�����;�����]�������������������̋�U��Q�E�    �tjP�ܑ�E��MQ���tj�E���]��������������̋�U��tjP�ܑ]��������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̋�U��E��w$���A���F���tRP�EQP�D   ��]útCR�   P�E�   QP�$   ��]�������������������������������̋�U���@  ��A3ŉE��ES�]VW�}S������������ǅ����    ��������������uS�d������������5�j j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ�����Gh  ��  ����������t%���������FPSQW�}  �����"  2��������� ������u���  ��t������   h  ������R������Ph  ������Q���S�J�������t-������������RWh�G������P�EQ������RP���   �=�j j h
  ������Qj�������Rj h��  ��G�ׅ�t������j j h
  ������Pj�������Qj h��  �xG�ׅ�t������������������������R�UPhPGVQSR����������u̋M�_^3�[�6�����]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�+h�d�    P��$SVW��A1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@����	�   Ëe��E������E�M�d�    Y_^[��]��������������������������������������̋�U��j�h�+h�d�    P��$SVW��A1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@����	�   Ëe��E������E�M�d�    Y_^[��]����������������������������������������������������̋�U���  ��A3ŉE��=�A��E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ���F������A��u�Њ@��u�W������+�O�OG��u��������ȃ���F�Ȋ@��u�������+���O�OG��u������ȃ��_��|H��A������SjPQ�������^[�M�3��+�����]��������������������������������������������������������������������̋�U���D  ��A3ŉE�S��AV�uW�}�����������   h�I� �����   h�IP����`]����   ����   �M�Vh�IQh�I��$Rh�I�~ Wh�Ih8I������hIQ�ЋV��$RW�E�P�M�Q��   ��8hI�U�RhI�E�PhI������Q���������R�`]������������PjSQ������(_^[�M�3��֡����]�h�HjSW�������M�_^3�[贡����]�����������������������������������������������������������������������������̋�U����ESV�u�E��EW3�+ƉE����M��r�   ;�s&�0�U���QhJR�`]�E��E����GF�ɋM�E�y� � _^[��]���������������������������������̋�U���  ��A3ŉE��=�A��E��   SV����   �ȍq�A��u�+΃�:��   ww������3Ɋ��F������A��u�Њ@��u�W������+�O�OG��u��������ȃ��G�Ȋ@��u�������+���O�OG��u������ȃ��_��J��ASjP�EP������^[�M�3�������]�����������������������������������������������������������������������̸   ����������̋�U��E��w	��(K]�3�]������̋�U��M��w�U���A���A]Ã��]�����������̋�U��M�d]�d]�h]    ]�����������������̋�U��M�h]�h]�d]    ]�����������������̡d]����������̡h]�����������u�U��� PRSVWh�Kh�KjBh@Kj�_�������u�_^[ZX��]������������������������̋�U�층�]����̋�U���]����̋�U��j jhHMhMh�Lh   h   j ������P�ί����]�������������������������̋�U��} u��EP�MQ�UR�EP�MQ胶��]������������������������̋�U��j �EP�޸����]�����������̋�U����EP�M��o����M�R輴������et�E���E�M�R�٢������u�E�Q茴������xu	�U���U�E��M��M�葢������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M��:�����]������������������������������������������������̋�U��Q�M��E��@ �} ��   貫���M��A�U��B�M��Pl��E��H�U��Ah�B�M��;LKt�E��H�Qp#�Hu
胲���M���U��B;�Ft�M��Q�Bp#�Hu�ƴ���M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������������������������������������������������������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]�������������������̋�U��Q�M��E���]����������������̋�U��j �EP������]�����������̋�U���V�EP�M������M���t*�E�0�M��U�������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��ğ������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M��n���^��]�������������������������������������������������������������������̋�U��Q�E�������Az	�E�   ��E�    �E���]���������������������̋�U����} t$�EP�MQ�U�R�Ԣ�����E�M���U��P��EP�MQ�U�R�D������E�M���]������������������������������̋�U��j �EP�MQ�UR�η����]�������������������̋�U���D��A3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�P�����3Ƀ} ���Mă}� u!h�Nj h�  hNj肞������u̃}� u3�����    j h�  hNh�Mh�N�]������   �  3�;E��ىM�u!h�Mj h�  hNj��������u̃}� u3諷���    j h�  hNh�Mh�M��������   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�������Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3��;�����]��������������������������������������������������������������������������������������������������������������������̋�U���@�E�    �E P�M�舧��3Ƀ} ���M܃}� u!h�Nj h3  hNj�x�������u̃}� u@�	����    j h3  hNhPh�N�S������E�   �M�芶���E���  3�;E��ىM�u!h�Mj h4  hNj��������u̃}� u@蔵���    j h4  hNhPh�M�ޮ�����E�   �M������E��}  3��} ����#E��	;E��ىM�u!h�Oj h<  hNj�~�������u̃}� u@����� "   j h<  hNhPh�O�Y������E�"   �M�萵���E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�V  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��&�������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  hNhPh�Nh�N�U�R�E�P�1�����P� ������M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE����j��t �U����0uj�M��Q�U�R�������E�    �M�蓳���Eċ�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�?�����]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M�葢���} }�E    3Ƀ} ���M��}� u!h�Nj h�  hNj�t�������u̃}� u@�����    j h�  hNh�Ph�N�O������E�   �M�膱���E���  3�;E��ىM�u!h�Mj h�  hNj���������u̃}� u@萰���    j h�  hNh�Ph�M�ک�����E�   �M������E��g  �E�  �M��;M��ډU�u!h0Pj h�  hNj耖������u̃}� u@����� "   j h�  hNh�Ph0P�[������E�"   �M�蒰���E���  �M��Q�4����%�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ�O������E��}� t�U� �E��E��M������E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ还�����E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M��r����E���  �M��Q�?��������� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4脮��%�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M��>�������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U������E�U��E܅���   �} ~}�M��Q���� #E�#U��M��@���f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U�������E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M�跬��f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4�ȫ��%�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R豑������0�M��U���Uj h�  �E�P�M�Q�9����E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�\����Ѓ�0�E��M���Mj jd�U�R�E�P�����E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�
����ȃ�0�U�
�E���Ej j
�M�Q�U�R蕐���E��U��E���0�M��U���U�E�  �E�    �M�襪���E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ腅����]���������̋�U��j �EP�MQ�UR�EP�MQ�Ņ����]�����������̋�U���D��A3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�`�����3Ƀ} ���Mă}� u!h�Nj h*  hNj蒍������u̃}� u3�#����    j h*  hNh�Ph�N�m������   ��   3�;E��ىM�u!h�Mj h+  hNj�*�������u̃}� u3軦���    j h+  hNh�Ph�M�������   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�?������Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�   ���EȋEȋM�3��b�����]�����������������������������������������������������������������������������������������������������������̋�U���4�E�H���M��UR�M�賖��3��} ���E�}� u!h�Nj h�  hNj裋������u̃}� u@�4����    j h�  hNh�Ph�N�~������E�   �M�赥���E��  3�;U��؉E�u!h�Mj h�  hNj�.�������u̃}� u@迤���    j h�  hNh�Ph�M�	������E�   �M��@����E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P��  ���M��0�U����U���E�M�H�M��} ��   j�U�R�  ���M�蔉��� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�  ���EPj0�M�Q�a������E�    �M�������EЋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�c�����]���������������̋�U���P��A3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�,�����3Ƀ} ���M��}� u!h�Nj ho  hNj�^�������u̃}� u3�����    j ho  hNh�Ph�N�9������   �i  3�;E��ىM�u!h�Mj hp  hNj���������u̃}� u3臡���    j hp  hNh�Ph�M�њ�����   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�������E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�?������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ��������M�3�诀����]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�A�����]�����������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�}�����E��{�}fu!�E P�MQ�UR�EP�MQ�������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�}�����E��#�U R�EP�MQ�UR�EP�MQ�~������E��E���]������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR�C~����]�����������������������̋�U��} t#�EP��������P�MQ�UUR�A�����]����������������̋�U��Q�E�    �	�E����E��}�
s�M����AR���M����A�ԋ�]�����������������̋�U��j
�����3�]����������̋�U��j�h ,h�d�    P���SVW��A1E�3�P�E�d�    j�������E�    �E�x ��   �t]�M��E�p]��U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�E������/�M�M��U�z uh�Qj jXh�Pj�D�������u�랋M�QR�������E�@    �E������   �j�ޑ����ËM�d�    Y_^[��]������������������������������������������������������������������������̋�U��j�h ,h�d�    P���SVW��A1E�3�P�E�d�    �E�x �L  h (  h�h��j �M��	Qj 膌�����E�}� u3��   �U�R訅�����E��E��M����M���v�U�U���� u�M�M�� ��j�G������E�    �U�z ��   j�Y������E܃}� ��   �E���P�=������E؋M�U؉Q�}� t[j h�   h�PhxRh�Q�E�P�M���Q�U�BP�\�����P�+������M܋U�B��M܋U�B�A�M�U܉Q��E�P�"������M�Q�l������E������   �j�������ËU�B�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������̋�U��j�h@,h�d�    P���SVW��A1E�3�P�E�d�    j讁�����E�    �E�x ��   �t]�M��E�p]��U��U�}� tY�E�M�;Qu�E��M�Q�P�E�P�;������2�M�M��U�z u!h�Qj h�   h�Pj��������u�뛋M�QR��������E�@    �E������   �j�{�����ËM�d�    Y_^[��]���������������������������������������������������������������������̋�U���E��u	� (  f�M�URh�h���EP�MQ�UR�N�����]���������������������̋�U��j�h`,h�d�    P���SVW��A1E�3�P�E�d�    �E�x �a  j�������E�    �M�y �*  h (  j �U��	Rj ��x�����E�}� u"�E�    j��E�Ph�A�������E��  �M�Q�Ɂ�����E��U��E����E���v�M�M���� u�E�E��  ��j�|�����E܃}� ��   �E�    �M���Q�|�����E؃}� taj h4  h�Ph,Sh�R�U�R�E���P�M�Q蠘����P�o������U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P賋�����M�Q觋�����E������   �j�4�����ËU�B�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������̋�U��j�h�,h�d�    P���SVW��A1E�3�P�E�d�    j��}�����E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P膊�����M�Q�z��������E������   �j������ËM�d�    Y_^[��]�����������������������������������������������̋�U��j ��]�����������������̋�U����]� ����������������̋�U��EP��AQ����]� �������������������̋�U���A]����̋�U��Q��AP���E��}� u ��]Q�ܑ�E��U�R��AP���E���]������������������������������̋�U��EP�MQ��]R�ܑ��]� ���������������̋�U���h�S���E��}� u跄��3���  h�S�E�P����|]h�S�M�Q�����]h�S�U�R�����]h�S�E�P�����]�=|] t�=�] t�=�] t	�=�] u,�|]2�����]����]����]����A�=�A�t��]Q��AR����u3���   �~~���|]P���|]��]Q����]��]R����]��]P����]�L�����u脃��3��   hr��|]Q�ܑ�У�A�=�A�u	�V���3��rh  hxSjh  j�������E��}� t�U�R��AP��]Q�ܑ�Ѕ�u	����3��(j �U�R�ȏ�����ؑ�M���U��B�����   ��]������������������������������������������������������������������������������������������������������������������������������������̋�U��=�A�t��AP��]Q�ܑ����A�����=�A�t��AR����A�����/r��]����������������������������̋�U��j�h�,h�d�    P���SVW��A1E�3�P�E�d�    h�S���E�E�@\`m�M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@hhBj�x�����E�    �M�QhR���E������   �j�������j�sx�����E�   �E�M�Hl�U�zl u�E�LK�Hl�U�BlP蚋�����E������   �j谅����ËM�d�    Y_^[��]��������������������������������������������������������������������������̋�U����$��E���AP�n���ЉE��}� u}j h�  hxSjh  j�5x�����E��}� tW�M�Q��AR��]P�ܑ�Ѕ�t%j �M�Q�Ό�����ؑ�U���E��@�����j�M�Q�V������E�    �U�R� ��E���]�����������������������������������������������������������̋�U��Q��p���E��}� u
j螊�����E���]�����������̋�U��j�h�,h�d�    P���SVW��A1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P�w������M܃y, tj�U܋B,P�]������M܃y4 tj�U܋B4P�C������M܃y< tj�U܋B<P�)������M܃y@ tj�U܋B@P�������M܃yD tj�U܋BDP��������M܃yH tj�U܋BHP�ۃ�����M܁y\`mtj�U܋B\P较����j�u�����E�    �M܋Qh�U��}� t%�E�P�(���u�}�hBtj�M�Q�y������E������   �j��������j�-u�����E�   �U܋Bl�E�}� t4�M�Q�3������U�;LKt�}�HJt�E�8 u�M�Q�o�����E������   �j�T������j�U�R�������M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��=�A�tO�} u)��AP����t��AQ��AR���ЉEj ��AP��]Q�ܑ�ЋUR��~���=�A�tj ��AP��]������������������������������������������̋�U���ؑ]���̋�U���,�]���̋�U��Q�EP�MQ�UR�@_P�MQ�,������E��E���]������������������̋�U��j j j�EP�MQ�������]�������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�D   ���E��}� u�}� t�������t
������M���E���]������������������������̋�U��Q�EP�MQ�UR�EP�MQ�   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP��~������u�} t	�M�   3��뗋�]�����������������������������̋�U��j j j�EP��{����]�������̋�U��j�h -h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    j�q�����E�    �=�] vU��]��9�]u6�xj����u!h�Uj h  hUj��o������u���]    ���]����]��A�E؃= B�t�M�; Bu̃=�N tu�UR�EP�M�Q�UR�EPj j��N����uP�} t%�MQ�URh�Tj j j j �+p������u�� h�Th@j j j j �	p������u��D  �U����  ��t��A��u�E�   �}�v3�MQh�Tj j j j��o������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t hHTh@j j j j�do������u̋M��$�MԋU�R�h�����E܃}� u�} t	�E�    �r  ��A����A�}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+�];Mv��]U��]�
��]������]E��]��];�]v��]��]�=�] t��]�M܉H�	�U܉�]�E܋�]��U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉�]j�BR�E܃�P��m����j�BQ�U�E܍L Q��m�����UR�BP�M܃� Q�m�����U܃� �U��E������   �j�{����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�(������E��}� u�}� t�3�����t
�*����U���E���]����������������������������̋�U��Q�} v�����3��u;Es�����    3��K�E�E�E�MQ�UR�EP�MQ�@_R�EP��������E��}� t�MQj �U�R�k�����E���]���������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�l�����E��}� u�}� t������t
�����M���E���]������������������������̋�U��Qj j j�EP�MQ�UR�Ha�����E��E���]����������������������̋�U��j�h -h�d�    P���SVW��A1E�3�P�E�d�    j�k�����E�    j�EP�MQ�UR�EP�MQ�b   ���E��E������   �j�gx����ËE�M�d�    Y_^[��]����������������������������������������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�Yb�����  �} t�}� u�EP�MQ�mx����3��  �=�] vV��]��9�]u6�;c����u!h�Uj h�  hUj�h������u���]    ���]����]��A�U�= B�t�E�; Bu̃=�N ty�MQ�UR�E�P�MQ�U�R�EPj��N����uR�} t%�MQ�URh,Yj j j j ��h������u�� h Yh@j j j j ��h������u�3��  �}��v`�} t)�UR�EP�M�Qh�Xj j j j�h���� ��u���E�Ph�Tj j j j�nh������u��=����    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URhPXj j j j�h������u�� hHTh@j j j j��g������u��Qj�BR�E�����P�  ����t1�MQh�Wj j j j�g������u��~����    3��t  �EP��h������u!h�Wj h  hUj�f������u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h�Vj h#  hUj�Of������u��d�M�Q����  ��u�E%��  ��u�E   �M��];Qs1�EPh�Vj j j j��f������u�����    3��  �} t%�U���$R�E�P�Th�����E��}� u3��_  �#�M���$Q�U�R�a�����E��}� u3��:  3�u���A����A�}� u|�=�]�s9�U�]+B��]���+�];M�v��]U���]�
��]�����E���]+H��]��]U���]��];�]v��]��]�U��� �U�E��M�;Hv$�U��E�+BP�BQ�U��E�BP�we����j�BQ�U�U�R�^e�����}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!h8Vj h�  hUj�Vd������u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8��];M�t!h�Uj h�  hUj��c������u̋E��H��]�U��z t�E��H�U����7��];M�t!h�Uj h�  hUj�c������u̋E����]�=�] t��]�E��B�	�M���]�U�]��M��A    �U���]�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es�;{���    3��g�E�E�E��} t�MQ�"l�����E��UR�EP�MQ�U�R�EP�v�����E�}� t �M�;M�s�U�+U�Rj �E�E�P��a�����E��]����������������������������������������������������̋�U��Qj j j�EP�MQ�}v�����E��E���]����������̋�U��j�h@-h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E��}� u!h�Yj h�  hUj�a`������u̃}� u-��y���    j h�  hUhpYh�Y�<s����3��c�}�v�y���    3��Nj�Sa�����E�    j �UR�EP�MQ�UR�EP�������E��E������   �j�n����ËE�M�d�    Y_^[��]�������������������������������������������������������������������̋�U��j�EP�rh����]�����������̋�U��j�h`-h�d�    P��SVW��A1E�3�P�E�d�    j�^`�����E�    �EP�MQ�h�����E������   �j�m����ËM�d�    Y_^[��]����������������������������������̋�U��Q�=�] vU��]��9�]u6��X����u!h�Uj h  hUj�m^������u���]    ���]����]�} u�l  �}uOj�BP�M�����Q�	  ����t/�URh`^j j j j��^������u��w���    �  �=�N tDj j j �MQj �URj��N����u%h@^h@j j j j �r^������u���  �MQ�_������u!h�Wj h*  hUj�t]������u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!h�]j h0  hUj�]������u̋�A���m  j�BP�M���Q�k  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��0TPh]j j j j�Z]����(��u��<�U��� R�E��HQ�U��B%��  ��0TQhh\j j j j�]���� ��u�j�BP�M��Q�E��L Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��0TPh�[j j j j�\����(��u��<�U��� R�E��HQ�U��B%��  ��0TQh [j j j j�b\���� ��u̋E��xue�M��y����u	�U��z t!hhZj hi  hUj�[[������u̋M��Q��$R�BP�M�Q��[�����U�R�Yi�����Q  �E��xu�}u�E   �M��Q;Ut!h Zj hw  hUj��Z������u̋M���]+Q��]��A����   �M��9 t�U���M��Q�P�6��];E�t!h�Yj h�  hUj�Z������u̋U��B��]�M��y t�U��B�M����5��];E�t!h�Yj h�  hUj�9Z������u̋U����]�M��Q��$R�BP�M�Q�Z�����U�R�-h�����(�E��@    �M��QR�BP�M��� Q�Z������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�EP�]����]�����������̋�U��j�h�-h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E܃}� u!h�Yj h�  hUj�X������u̃}� u1�q���    j h�  hUh�^h�Y��j��������8  �=�] vV��]��9�]u6�R����u!h�Uj h�  hUj�W������u���]    ���]����]j�X�����E�    �UR�jY������u!h�Wj h�  hUj�9W������u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!h�]j h�  hUj��V������u̋E��xu�}u�E   �M��Q�U��E������   �j�se����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������̋�U��Q� B�E��M� B�E���]������������������̋�U��j�h�-h�d�    P���SVW��A1E�3�P�E�d�    j��V�����E�    �EP�W������te�M�� �M�U�B%��  ��tC�M�yt:�U�B%��  ��t*�M�yt!h�]j h?  hUj�7U������u̋E�M�H�E������   �j��c����ËM�d�    Y_^[��]�������������������������������������������������������������̋�U��Q��N�E��M��N�E���]������������������̋�U�졀N]����̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�����������������������̋�U��j�h�-h�d�    P���SVW��A1E�3�P�E�d�    ��A��u
�   ��  j�*U�����E�    �LV���E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$�Yh|ah@j j j j �HT������u��   hPah@j j j j �#T������u��dh(ah@j j j j �T������u��Bh ah@j j j j ��S������u�� h�`h@j j j j �S������u��E�    ��  �E�   ��]�E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��0T�U���E��`j�BP�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh]j j j j ��R����(��u��-�E�� P�M�QR�E�Phh\j j j j �R���� ��u��E�    j�BR�E�H�U�D
 P�2�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph�[j j j j �5R����(��u��-�U�� R�E�HQ�U�Rh [j j j j �R���� ��u��E�    �M�y ��   �U�BP�BQ�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� Rh `j j j j �Q���� ��u��"�M�� Qh`_j j j j �sQ������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rh_j j j j �"Q����(��u��-�M�QR�E�� P�M�Qh�^j j j j ��P���� ��u��E�    �G����E������   �j��^����ËE܋M�d�    Y_^[��]ÍI �U�U{UVU���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�-h�d�    P���SVW��A1E�3�P�E�d�    ��A�E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h�aj hy  hUj�;N������u̃}� u0��g���    j hy  hUh�ah�a�a������A�sj�?O�����E�    ��A�M�}�t7�U��t��]   ��E��%��  ��]��]    �M��A�E������   �j�c\����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��j�h .h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E��}� u!h�cj h�  hUj��L������u̃}� u+�Rf���    j h�  hUh�ch�c�_�����s��A��u�fj�M�����E�    ��]�E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j��Z����ËM�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��3��} ��]����������������̋�U��} u3��1j j �E�� P�4S������u3���M�� Qj �<_R�0�]������������������������������̋�U��j�h .h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP��L������u3���   j��K�����E�    �M�� �M��U��B%��  ��t"�M��yt�U��B%��  ��t	�M��yukj�UR�EP�R������tU�M��Q;UuJ�E��H;�A<�} t�U�E��H�
�} t�U�E��H�
�} t�U�E��H�
�E�   ��E�    �E������   �j�X����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U��Q�EP�`K������u�����M�� �M��U��B��]������������������̋�U��Q��]�E��M��]�E���]������������������̋�U�졤]]����̋�U��j�h@.h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E܃}� u!h�dj h�  hUj�H������u̃}� u.�b���    j h�  hUhldh�d�\[�����m  j�I�����E�    �U��]��E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡ�]�E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�Rh dj j j j ��G���� ��u���M�Qh�cj j j j ��G������u������E��]�H,�U��]�B0�E������   �j�U����ËM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E�}� u!h�dj h�  hUj�F������u̃}� u0�_���    j h�  hUheh�d��X����3��  3҃} �U��}� u!h�dj h�  hUj�E������u̃}� u0�+_���    j h�  hUheh�d�uX����3��0  3Ƀ} ���M�}� u!h�dj h�  hUj�1E������u̃}� u0��^���    j h�  hUheh�d�X����3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u��A��t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��hN���M���B��P�MQ�#   ���M��]����]��������������������̋�U��j�h`.h�d�    P���SVW��A1E�3�P�E�d�    �E�    j�WD�����E�    h0fh@j j j j �C������u̃} t�M��Uࡠ]�E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u��A��u��  �U�z twj j�E�HQ�J������tj�U�BP�4���t$�M�QRhfj j j j ��B������u��)�M�QR�E�HQhfj j j j �B������u̋E�HQh fj j j j �B������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph�ej j j j �OB���� ��u̃=�] t,j�U�� R�4���u�E�HQ�U�� R��]����E�P�MQ�  ���   �U�zu;�E�HQ�U�� Rh�ej j j j ��A������u̋M�Q�UR�x  ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� PhTej j j j �wA���� ��u̋U�R�EP�  ��������E������   �j�OO�����h8eh@j j j j �)A������u̋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���t��A3ŉE��EP�M��EJ���E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M��w>����t3�M��k>������   ~ �M��X>��PhW  �E�P�S�����E��hW  �M�Q�M��.>��P��7�����E��}� t	�U��U���E�    �E��M��L��=X����U��3X���     �E�PhJ�M�k��1   +�R�E�k��L�Q��M������}*j h	  hUhxfh\fj"j��W���R��9���� ��W���M��������U��D� �E�P�M�QhHfj j j j ��>������u̍M��FX���M�3���7����]������������������������������������������������������������������������������������������������������������������̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP��O���E]������������������̋�U���8��A3ŉE��E�P�pB�����}� u�}� u��A��t7�}� t1h�fh@j j j j �=������u�j �fP�����   �3��M�3��6����]������������������������������������̋�U���3��} ���E��}� u!h�dj h�	  hUj�K<������u̃}� u.��U���    j h�	  hUh8gh�d�&O�����   �E�    �	�U����U��}�}>�E���0TQ�U��E�L�Q�U��E�L�Qhgj j j j �<���� ��u�볋E�H,Qh�fj j j j �g<������u̋E�H0Qh�fj j j j �E<������u̋�]�������������������������������������������������������������������̋�U��j j j �EP�MQ�(<����]�������������������̋�U��EP�MQj �UR�EP��;����]���������������̋�U��j j j �EP�MQ�UR�t;����]���������������̋�U��j j j �EP�MQ�UR�EP�C����]�����������̋�U��EP�MQj �UR�EP�MQ�;����]�����������̋�U��EP�MQj �UR�EP�MQ�UR�$C����]�����������������������̋�U��j j �EP�MQ�UR��:����]�����������������̋�U���(�E��#E������E�u!h�gj h�
  hUj�9������u̃}� u0�)S���    j h�
  hUh�gh�g�sL����3��@  �} t�U;Ur	�E�    ��E�   �E܉E��}� u!hlgj h�
  hUj�9������u̃}� u0�R���    j h�
  hUh�ghlg��K����3��   �}v�U�U���E�   �E؃��E3�+M���M�U�E�L�M��UU��U�E;E�v�1R���    3��i�MQ�URj�E�P�1�����E�}� u3��F�M�M�M�U��#�+M�M��E�+E���E�j�BQ�U���R��8�����E��M��E���]������������������������������������������������������������������������������������������������������������������������̋�U��j j �EP�MQ�UR�EP�B8����]�������������̋�U��j j �EP�MQ�UR�EP�MQ�V@����]���������̋�U���4�} u!�EP�MQ�UR�EP�MQ�)8�����  �} u�UR�DQ����3��  �E������E�j�BQ�U��R�V�������t1�EPh�hj j j j�~7������u��MP���    3��C  j�BR�E���P��������u�MQhdhj j j j�07������u̋E��#E������E�u!h�gj h�  hUj�26������u̃}� u0��O���    j h�  hUh hh�g�I����3��  �} t�U;Ur	�E�    ��E�   �EԉE؃}� u!hlgj h�  hUj�5������u̃}� u0�BO���    j h�  hUh hhlg�H����3��  �U��P�@�����M��U++E�}v�E�E���E�   �MЃ��M3�+U���U�E�M�T�U�EE�E�M;M�v�N���    3��   �UR�EPj�M�Q�).�����E��}� u3��   �U�U�U�E��#�+U�U��M�+M���M�j�BR�E���P�O5�����M��U���E�;Ev�M�M���U�ŰE�P�MQ�U�R��>����j�E��Q��C�����E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es��L���    3��s�E�E�E��} t�MQ�UR�EP�G�����E��M Q�UR�EP�MQ�U�R�EP��3�����E�}� t �M�;M�s�U�+U�Rj �E�E�P�3�����E��]��������������������������������������������������������̋�U��EP��L����]�������������̋�U��Q�} u�   �E������E�j�BQ�U��R���������t!�EPhij j j j��2������u��Lj�BR�E���P��������u�MQhdhj j j j�2������u�j�E��Q�LA������]�����������������������������������������������������̋�U��Q��A�E��M��A�E���]������������������̋�U��Q��]�E��E���]�����������̋�U�졬]]����̋�U��EP�MQ�UR�L/����]���������������������̋�U��� �E�    �E�    �E�    �E�    �E�    3��} ���E�}� u!h�ij h�  hUj�0������u̃}� u.�IJ���    j h�  hUh\ih�i�C��������w�E�    �U������U��E��Q�;�����E��U��E+�E�3�+M���M�}v�U�U���E�   �E����E�M�U�D
+E�E�M�+M�+M�M��E���]�������������������������������������������������������������������̋�U��Q�=�B th�B�D������t�EP��B���=��h05h3�I�����E��}� t�E��Gh���/����h2h 0�R  ���=�� th���3D������tj jj ���3���]���������������������������������������������������̋�U��j j �EP�>  ��]���������̋�U��j j�EP�  ��]���������̋�U��jj j �   ��]�����������̋�U��jjj ��  ��]�����������̋�U���TB���EP�1����h�   �'1��]��������������̋�U��Q��]�E��	�M����M��}� t�U��: tj�E��Q�|=������j��]R�i=������]    ��]�E��	�M����M��}� t�U��: tj�E��Q�.=������j��]R�=������]    j��]P�=����j��]Q��<����j���R�ܑP��<������]    ��]    ��3�������FP�(���u'�=�FhBtj��FQ�<������FhB��FR����]�����������������������������������������������������������������������������������������������̋�U��j�h�.h�d�    P���SVW��A1E�3�P�E�d�    �P=���E�    �=�]�U  ��]   �E��]�} ��   ���Q�ܑ�E�}� ��   ���R�ܑ�E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�N2���U�9u��E�;E�s�h�M؋R�ܑ�E��'2���M؉�U܋��R�ܑ�EС��P�ܑ�E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���hH9h46�A  ��hP;hL:�/  ���=�] u#j��*������ t��]   �;$���9���E������   ��} t��$��Ã} t���]   ��$���MQ��-�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������̋�U���h�i���E��}� th�i�E�P����E��}� t�MQ�U���]�����������������̋�U��EP��$�����MQ�8�]�������������������̋�U��j��*����]���������������̋�U��j�T8����]���������������̋�U��Q��/���E��E�P�� �����M�Q�@�����U�R�43�����E�P�+!�����M�Q��+�����U�R��2������]����������������������̋�U��E;Es�M�9 t�U��ЋM���M��]�����������������������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�����������������̋�U���3��} ���E��}� u!h�jj h�  h0jj�;(������u̃}� u0��A���    j h�  h0jhjh�j�;�����   �y3҃=�] �U��}� u!h�ij h�  h0jj��'������u̃}� u0�`A���    j h�  h0jhjh�i�:�����   ��M��]�3���]������������������������������������������������������������������̋�U���3��} ���E��}� u!h�jj h�  h0jj�'������u̃}� u0�@���    j h�  h0jh�jh�j��9�����   �y3҃=�] �U��}� u!h�jj h�  h0jj�&������u̃}� u0�0@���    j h�  h0jh�jh�j�z9�����   ��M��]�3���]������������������������������������������������������������������̋�U���p�E�P�L�h�   hkjj@j ��>�����E��}� u�����  �M�����<�    �	�U���@�U����   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M��<�;U���   h�   hkjj@j �=�����E��}� u�<��E��   �M��U������<��� �<��	�M���@�M��U�����   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R�H���t[�E����M���������M��U��E���
�U��E���Jh�  �U���R�D���u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M������M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P�@��E��}����   �}� ��   �M�Q�H��E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�D���u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A������<�R�<�3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �	�E����E��}�@}y�M��<��� tg�U������E��	�M���@�M��U�����   9E�s�M��y t�U���R�P���j�E�����Q��/�����U�����    �x�����]���������������������������������������������������̋�U����=�� u����E�    �L]�E��}� u����e  �M����t,�E����=t	�U����U��E�P�8#�����M��T�U���juh ljj�E���P�z8�����E�M��]�=�] u�����   �L]�U��	�E�E��E��M������   �E�P��"�������E��M����=��   j~h ljj�E�P�8�����M��U�: uj��]P�|.������]    ����rj h�   h�kh�khLk�M�Q�U�R�E�Q�9����P�x*�����U���U��B���j�L]P�.�����L]    �M��    ���   3���]��������������������������������������������������������������������������������������������������������������������̋�U����E�    �=�� u����_ h  h ^j �T�h ^������=�� t������t����U���E� ^�E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   h\lj�M��U���P������E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�   ���U�����]�E���]3���]�������������������������������������������������������������������������̋�U��E��]]�����������������̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�*������t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P�(������t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R�Q(������t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �\��E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j ���E��}� tjJh�lj�M�Q�������E�}� u�U�R�X�3��Dj j �E�P�M�Q�U�R�E�Pj j ����uj�M�Q��&�����E�    �U�R�X��E��]������������������������������������������������������������������������̋�V��$��=�&s���t�Ѓ����&r�^����������̋�V� (��=\*s���t�Ѓ���\*r�^����������̋�U��Q�E�   j h   j �`��<_�=<_ u3���   ��]�������������������������̋�U��<_P�d��<_    ]�������������������̋�U��=<_ uhHmj jhh�lj�
������u̡<_]�������������̋�U���0�E� �E�   �E���E��M����M�U��B3�A�EԋM�Q�U�R��  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M��s���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=8 t h8��)������tj�UR�8���M����U��*���E��H;M�th�A�U�R�M����U�����E��M�H�U�R�E�P��   ���U�M�I�t�������&�U��z�th�A�E�P�M������������E��M߅�t�U�R�E�P�   ���E��]������������������������������������������������������������������������������������������������������������������������̋�U����E�8�t%�M��E��M��U�EB3E��E��M�����M�Q�E��M��U�EB3E��E��M��h����]���������������������������������̋�U����E�    �E�    �=�AN�@�t��A%  ��t��A�щ�A�   �U�R�t��E��E�M�3M��M��p�3E�E��ؑ3E�E��l�3E�E�U�R�h��E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M��A�U��҉�A��]����������������������������������������������������������������̋�U��}csm�u�EP�MQ�o'������3�]����������̋�U����!���E��}� u3���  �E��H\Q�UR�S  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  ��m�U��	�E����E���m�m9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��;Ut�E����E���mk�M9M�s�ڋ�mk�U9U�s
�E��;Mt3���E���]�������������������������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������������������������������������������������������̋�U���(  �P`�L`�H`�D`�5@`�=<`f�h`f�\`f�8`f�4`f�%0`f�-,`��``�E �T`�E�X`�E�d`��������_  �X`�T_�H_	 ��L_   ��A��������A����������_j�7����j ���h n����=�_ u
j�����h	 ��|�P�x���]����������������������������������������������������������������������������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uhoj jph�nj�Z������u̃}� u.��%���    j jph�nh�nho�8��������)  �} t�} u	�E�    ��E�   �M̉MЃ}� uh0nj jsh�nj��������u̃}� u.�q%���    j jsh�nh�nh0n���������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R������E��} u�E��P�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �g�����EċE���]�������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�	!����]���������������̋�U��Q�E�    �\B��t
j
������4���E��}� t
j�������\B��tjh  @j� ����j������]��������������������������������̋�U��Q�\B�E��M��#M��U#Uʉ\B�E���]���������������������̋�U��j�������tj�������u#�=X]uh�   �����h�   �����]�������������������������̋�U��Q�E�    �	�E����E��}�s�M��U;�Xyu�E���\y���3���]�������������������������������̋�U���   ��A3ŉE�EP������E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j�o���������������� t������t���E�   ��E�   �}� ��  j�V������tj�G��������   �=X]��   j��@��E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P�����P������Q�U�R�����  �}�   ��  ǅ����Bc������-c���  +ȉ�����������������j h  hh~hH~hx}h4}h  hc�!����P������3�������f��  h  ������Rj �����u:j h  hh~hH~h�|hh|������P������Q�J!����P�d����������R�	��������<vk������P�	�����������TA�������j h  hh~hH~h�{jh�{������+�������������+�Q������R�l����P������j h  hh~hH~h0{h({h  hc�=�����P�����j h  hh~hH~h�z�E�Ph  hc������P�w����h  h0zhc�g �����M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   ��A3ŉE�}��  �E�E���p����M�ǅd���    ǅh����   ��h���R�E�P�MQ�UR�EP��������l�����l��� ��   �$���zt�  j j �MQ�UR�EP�D�������h�����h��� u��   j^h�jj��h���Q�������E��}� u��   ǅd���   ��h���R�E�P�MQ�UR�EP���������l�����l��� u�   jih�jj��l���Q�~�����U���E��8 u�]j jlh�hdh�~��l�����Q�U�R��l���P�M��R�� ����P�������d��� tj�E�P�����3��-  ��d��� tj�M�Q���������  �  �}��   �U��\�����\����     j j �MQ�UR�����`�����`��� u�Zh�   h�jj��`���P�������\������\����: u�(��`���P��\����R�EP�MQ�����u�3��mj��\����P��������\����    ����I�D�} u>ǅX���    j��X���R�E    P�MQ�����u�����U��X����3������M�3�������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�tj]�����������������̋�U��E�U��DV�u�     j�E�P3�NVf�
�����u3�^��]ËM�U�E�QRP�����t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=|j u �=xj uH�  �xj��t:�|j��xjh��P���3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�Rh��V�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ���P��������   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ���P����M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ��A3ŉE��=}j t3��M�3�������]��}j��   ����   VWh`����= ��5����t?h  ������QP�օ�t,h  ������R������P��  ����t������Q�ׅ�uBh  ������Rj �օ�t,h  ������P������Q�  ����t������R�ׅ�u3�_^�M�3��������]����������������������������������������������������������������̋�U���  ��A3ŉE�Vh|�� �����u^�M�3��Q�����]�W�=��hl�V�׉�������u_^�M�3��(�����]�ShX�V�׋؅�t4hH�V�׋���t&������Pjj h؀h  ���������tV���[_3�^�M�3��������]Í�����Q������������R������Pj h��Qǅ����  �Ӌ�����R����V�����u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M����D��H���E������L��H�P��P�T��H�X��Pf�\��Hf�P������P� ��M�[_3�^�������]����������������������������������������������������������������������������������������������������������������������̋�U���  ��A3ŉE��EV�uh   ������Qh   ������Rh   ������Qj�U�RP�|�����$��t3�^�M�3��������]�h��������j	P�f������u�h��������jQ�L������u�������R������P�E������Q�U�RPV����M������3�@^������]��������������������������������������������������������������̋�U��j�h�.h�d�    P���SVW��A1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh��j jah�j���������u̃}� u.�_���    j jah�hԂh�����������h  3҃} �U؃}� uh��j jbh�j�j�������u̃}� u.�����    j jbh�hԂh���H��������  j�p������E�    �,��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�,�j�U�R�������43�uh8�j jh�j�_�������u��E����������    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;,�tM�U�z t�E�H�U���M��E�H�J�U��    �E�,��H�,��E��M�,��h�   h��jj��������E�}� u�E������>���    �L�U��    �E�,��H�=,� t�,��E��M��A   �E�   �U�E�B�M�,��E������   �j�����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�	������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR�I����]���������̋�U��P  ������A3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �T���u8j h<  h�h��h��hd�h  ������Q�&����P��������������U��E�P��������@v]�M�Q�������U��D��E�j hE  h�h��hX�j�`BQ�U�������+й  +�Q�U�R� ����P�~������} t'�EP�.�������@v�MQ�������U�DÉE��;����������.���     �}uǅ����ȅ�
ǅ�����K�U���t�M�������
ǅ�����K�U���t�}uǅ�������
ǅ�����K�M���tǅ�������
ǅ�����K�} t�E�������
ǅ�����K�} tǅ�������
ǅ�����K�} t�M�������
ǅ�����K�} tǅ�������
ǅ�����K�}� t�U��������'�} t�E�������
ǅ�����K�������������}� tǅ�������
ǅ�����K�} tǅ�������
ǅ�����K������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U���Ph(�h�  h   ������Q������D�E�}� }*j h`  h�h��h\fj"j�'���R������ �����������}� }8j he  h�h��hp�h<�h   ������R�����P�������h  h�������P�������������������uj�������j�����������u�   �3��M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�.h�d�    P���SVW��A1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uh��j jah�j�^�������u̃}� u.�����    j jah�h��h���<��������h  3҃} �U؃}� uh��j jbh�j���������u̃}� u.����    j jbh�h��h������������  j� ������E�    �(��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�(�j�U�R�������43�uh8�j jh�j���������u��E���������    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;(�tM�U�z t�E�H�U���M��E�H�J�U��    �E�(��H�(��E��M�(��h�   h��jj�������E�}� u�E����������    �L�U��    �E�(��H�=(� t�(��E��M��A   �E�   �U�E�B�M�(��E������   �j������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP��������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR������]���������̋�U��X"  �"�����A3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj �����u8j h<  h�h�hx�hh|h  ������R�i����P�������������E��M�Q���������@v`�U�R�������M��TA��U�j hE  h�h�hX�j�dBP�M�������+����  +���P�M�Q�>�����P�	������} t'�UR�U�������@v�EP�D������M�TA��U������ ����������     �}uǅ����`��
ǅ����\��M���t�E�������
ǅ����\��M���t�}uǅ����<��
ǅ����\��E���tǅ����({�
ǅ����\��} t�U�������
ǅ����\��} tǅ����(��
ǅ����\��} t�E�������
ǅ����\��} tǅ������
ǅ����\��}� t�M��������'�} t�U�������
ǅ����\��������������}� tǅ�����{�
ǅ����\��} tǅ�������
ǅ����\�������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M��x�Rh0�h�  h   ������P�c�����D�E�}� }*j h`  h�h�h\fj"j����Q������ �����������}� }8j hc  h�h�hx�h�h   ������P�S����P�m�����h  h��������Q�[�����������������uj�L�����j�X���������u�   �3��M�3��h�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�d������E��E�    �E���]�����������������̋�U����E%�����E�M#M��������   �} tj j �k������U�3�t	�E�   ��E�    �M��M��}� uh؍j j1hH�j��������u̃}� u-�-����    j j1hH�h$�h؍�z������   �/�} t�EP�MQ��������U���EP�MQ�������3���]����������������������������������������������������������������̋�U��E��j]�����������������̋�U��Q��j�E��M�Q�ܑ�E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�#�����]����������������������̋�U��jh �j�a�����h ��|�P�x�]����������������������̋�U���8  ��A3ŉE��}�t�EP�������ǅ����    jLj ������Q�������������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M���������E�j ����U�R������������� u�}� u�}�t�EP��������M�3��������]�������������������������������������������������������������������������������������������������̋�U��Q�E�    ��j�E��M�Q�ܑ�E��UR���E�E��j�E���]������������������̋�U��Q�E�    ��j�E��M�Q�ܑ�E��E���]�����������������������̋�U��EP�MQ�UR�EP�MQ�������]�������������̋�U��EP�MQ�UR�EP�MQ�;���]����������������̋�U����EP�M��O����M��������t2�M���������   ~�M�����Ph  �UR��������E��h  �EP�M�����P�/������E�M�M�M��Y����E��]��������������������������������������������̋�U��=�m uh  �EP�A�������j �MQ�!�����]�������������̋�U����EP�M��_����M��������t/�M����������   ~�M�����Pj�UR��������E��j�EP�M�����P�E������E�M�M�M��o����E��]����������������������������������̋�U��=�m uj�EP�d�������j �MQ�������]����������������̋�U����EP�M������M��������t/�M����������   ~�M������Pj�UR�������E��j�EP�M�����P�e������E�M�M�M������E��]����������������������������������̋�U��=�m uj�EP��������j �MQ�������]����������������̋�U����EP�M������M�������t/�M��
�������   ~�M������Pj�UR�&������E��j�EP�M������P�������E�M�M�M������E��]����������������������������������̋�U��=�m uj�EP��������j �MQ�������]����������������̋�U����EP�M������M��6�����t2�M��*�������   ~�M�����Ph�   �UR�C������E��h�   �EP�M������P�������E�M�M�M�������E��]��������������������������������������������̋�U��=�m uh�   �EP��������j �MQ� �����]�������������̋�U����EP�M�������M��F�����t/�M��:�������   ~�M��'���Pj�UR�V������E��j�EP�M�����P�������E�M�M�M�������E��]����������������������������������̋�U��=�m uj�EP���������j �MQ������]����������������̋�U����EP�M�������M��f�����t/�M��Z�������   ~�M��G���Pj�UR�v������E��j�EP�M��%���P��������E�M�M�M�������E��]����������������������������������̋�U��=�m uj�EP���������j �MQ������]����������������̋�U����EP�M������M�������t2�M��z�������   ~�M��g���Ph  �UR�������E��h  �EP�M��?���P��������E�M�M�M������E��]��������������������������������������������̋�U��=�m uh  �EP��������j �MQ�������]�������������̋�U����EP�M������M�������t2�M���������   ~�M��w���PhW  �UR�������E��hW  �EP�M��O���P��������E�M�M�M��)����E��]��������������������������������������������̋�U��=�m uhW  �EP��������j �MQ������]�������������̋�U����EP�M��/����M�������t2�M���������   ~�M�����Ph  �UR�������E��h  �EP�M��_���P�������E�M�M�M��9����E��]��������������������������������������������̋�U��=�m uh  �EP�!�������j �MQ������]�������������̋�U����EP�M��?����M�������t/�M���������   ~�M�����Pj �UR��������E��j �EP�M��u���P�%������E�M�M�M��O����E��]����������������������������������̋�U��=�m uj �EP�D�������j �MQ�z�����]����������������̋�U��}�   ���]��������������̋�U��E��]���̋�U��Q�EP�MQ���������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP�n�������u�}_t	�E�    ��E�   �E���]�������������̋�U��Q�EP�MQ�U�������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP���������u�M��_t	�E�    ��E�   �E���]�������������������������̋�U��E�� ]���̋�U���4�EP�M�������}   ��   �M��Y�����t/�M��M�������   ~�M��:���Pj�UR�i������E��j�EP�M�����P��������Ẽ}� t,�M����������   �E��M��M�������E��*  ��U�U܍M�������E��  �M������ ���   ~D�M�����P�M�����   Q��������t"�U�����   �U��E�E��E� �E�   ������ *   �M�M��E� �E�   j�M��G�����BPj�M�Q�U�R�E�Ph   �M��&�����QR�M�����P������$�E�}� u�E�E؍M�������E��A�}�u�M��MԍM�������E��'��U��E���ЉUЍM������E���M�������]����������������������������������������������������������������������������������������������������������������������������̋�U��Q�=�m u$�}A|�}Z�E�� �E���M�M��E���j �UR���������]���������������������������̋�U��j�h�.h�d�    P���SVW��A1E�3�P�E�d�    �Z����E��E��Hp#�Ht�U��zl ��   j�[������E�    �E��Hh�M�U�;�FtI�}� t%�E�P�(���u�}�hBtj�M�Q�>������UࡐF�Bh��F�M�U�R���E������   �j�h�������	�E��Hh�M�}� u
j �������E�M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h /h�d�    P���SVW��A1E�3�P�E�d�    �E����������E��~����E܋Hh�M��UR��  ���E�E��M;H�  hN  h�jh   ��������E��}� ��  �U܋rh��   �}��E��     �M�Q�UR�I������E؃}� ��  �E܋HhQ�(���u�U܁zhhBtj�E܋HhQ�������U܋E��Bh�M܋QhR���E܋Hp���-  ��H���  j�5������E�    �E��H��j�U��B��j�M��Q��j�E�    �	�E���E�}�}�M�U�E�f�TPf�M�j���E�    �	�E���E�}�  }�M�M�U�A���D���E�    �	�M���M�}�   }�U�U�E䊊  ���E�׋�FR�(���u�=�FhBtj��FP�v������M���F�U�R���E������   �j��������(�}��u"�}�hBtj�E�P�+������U����    ��E�    �E؋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h8�
d�    P��$��A3�P�E�d�    �E�    �E�P�M������E�    ��j    �}�u)��j   ����E��E������M�������E��}�c�}�u)��j   ����E��E������M������E��N�4�}�u.��j   �M�������Q�U��E������M��^����E���E�E��E������M��D����EЋM�d�    Y��]����������������������������������������������������������������������������̋�U���,��A3ŉE�V�EP�������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0���F;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E���¨F�M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E����F�UU��B��MM��A����v����U�E�B�M�A   �U�BP��  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��p�Ff�DJ�ӋMQ�C  ��3��  �����} t!�}��  t�}��  t�UR�����u����k  �E�P�MQ������9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�\  ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=�j t�EP�  ��3�����^�M�3��R�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���  �M��}�w-�U������$����  ��  ��  �	�  �3���]ÍI ���������� ������������������������������������̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U����B�A���E�    �	�M����M��}�   }�UU��E����C��  �׋�]���������������������������������������������������������̋�U���(  ��A3ŉE�������P�M�QR������-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj ������ j �M�QRh   ������Ph   ������Qh   �U�BPj �������$j �M�QRh   ������Ph   ������Qh   �U�BPj ������$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3�苾����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��x����M�������H�y t �M�������P�B�E�M�������E����E�    �M������E���M�������]������������������������������������̋�U��=�� uj����������   3�]����������̋�U��Q�EP���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���E�    �	�M����M��}�m�U����E�|H�Ht$�M����U�|
P t�E����M�TPR���E����M�|L t$�U����E�|T t�M����U�D
TP��넋M���   �´   R����]���������������������������������������������������������������������������������̋�U��Q�} �  �EP�(��M���    t�U���   P�(��M���    t�U���   P�(��M���    t�U���   P�(��M���    t�U���   P�(��E�    �	�M����M��}�m�U����E�|H�Ht$�M����U�|
P t�E����M�TPR�(��E����M�|L t$�U����E�|T t�M����U�D
TP�(�넋M���   �´   R�(��E��]������������������������������������������������������������������������������������̋�U��Q�E���    ��   �M���   �N��   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P��������M���   R�������E���    t4�M���   �: u&j�E���   Q�������U���   P������j�M���   R������j�E���   Q�������U���    to�E���   �9 uaj�U���   -�   P�M�����j�M���   ��   R�3�����j�E���   ��   Q������j�U���   P�������M���   �Ht8�U���   ���    u&�M���   R�������j�E���   Q�������E�    �	�U����U��}���   �E����M�|H�Ht:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP�U������M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!hЎj h�   hX�j臽������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ�����������j�UR��������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR��������}� t�E�P�������}� t�M��9 u�}�HJt�U�R�׷�����E��]������������������������������������������̋�U��j�hP/h�d�    P���SVW��A1E�3�P�E�d�    �����E��E��Hp#�Ht	�U��zl uDj诼�����E�    �LKP�M���lQ�������E��E������   �j���������G����Pl�U�}� u
j �<������E�M�d�    Y_^[��]�����������������������������������������������������������̋�U���@��A3ŉE��E�    �E�    �EP�M��w����M�����Pj j j j �MQ�U�R�E�P� ����� �E��MQ�U�R�P������E��E���u8�}�u�E�   �M������E��j��}�u�E�   �M��v����E��N�:�M���t�E�   �M��X����E��0��U���t�E�   �M��:����E���E�    �M��&����E��M�3��Ƴ����]�������������������������������������������������������������������������������̋�U��j �EP�MQ迼����]�������̋�U���@��A3ŉE��E�    �E�    �EP�M������M��~���Pj j j j�MQ�U�R�E�P������ �E��MQ�U�R�������E��E���u8�}�u�E�   �M��"����E��j��}�u�E�   �M������E��N�:�M���t�E�   �M�������E��0��U���t�E�   �M�������E���E�    �M������E��M�3��V�����]�������������������������������������������������������������������������������̋�U��j �EP�MQ������]�������̋�U���@��A3ŉE��E�    �E�    �EP�M������M�����Pj j j j �MQ�U�R�E�P�@����� �E��MQ�U�R�������E��E���u8�}�u�E�   �M������E��j��}�u�E�   �M������E��N�:�M���t�E�   �M��x����E��0��U���t�E�   �M��Z����E���E�    �M��F����E��M�3�������]�������������������������������������������������������������������������������̋�U��j �EP�MQ�s�����]�������̋�U����E�E��M�Q�U�3��} ���E�}� uh�Nj j7hx�j�/�������u̃}� u0������    j j7hx�h\�h�N�������   �$  3�;U��؉E�uh�Mj j8hx�j�͵������u̃}� u0�^����    j j8hx�h\�h�M�������   ��  �U� 3��} ����#E��;E��ىM�uhؔj j=hx�j�U�������u̃}� u0������ "   j j=hx�h\�hؔ�3������"   �J  3��} ���E�}� uh��j j>hx�j��������u̃}� u0�����    j j>hx�h\�h����������   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R�]�������P�E��P�MQ落����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V�)����M��UR��������������0^]������������������������̋�U��Q�E�    �	�E����E��}�-s�M��U;�`Ku�E���dK�7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]��������������������������������������������̋�U��Q�s����E��}� u	�   ��������M�3���]�������������������̋�U��Q3��} ���E��}� u!h�jj h�   h�j�ͱ������u̃}� u%j h�   h�h�h�j�������   ��9����U� �3���]������������������������������������������̋�U��Q蓬���E��}� u	�   ���R����M�3���]�������������������̋�U��Q3��} ���E��}� u!h�jj h�   h�j��������u̃}� u%j h�   h�h��h�j��������   ��˷���U� �3���]������������������������������������������̋�U��Q賫���E��}� u	��L���E�����]���������̋�U��Q胫���E��}� u	��L���E�����]���������̋�U���,��A3ŉE��EP�M�Q�������U�Rj j���ċMԉ�U؉Pf�M�f�H�	������U�B�E�M��U��E�Pj j(h0�h�h���M�Q�UR�EP�q�����P�@������M�U�Q�E�M�3��z�����]���������������������������������������������������̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]����������������������������������������������������������������������������������������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�L�����   u������r)��$����Ǻ   ��r����$����$�����$�d���� �D�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l������$���I �Ǻ   ��r��+��$�p��$�l���������F#шG��������r�����$�l��I �F#шG�F���G������r�����$�l���F#шG�F�G�F���G�������V�������$�l��I  �(�0�8�@�H�P�c��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l���|��������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����j�E��M�����Ƀ��M�uhp�j j*h�j��������u̃}� u+�����    j j*h�h��hp���������E���E��j�E���]��������������������������������̋�U�졨j]����̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�j jh��j�X�������u̃}� u0������    j jh��ht�h��6������   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U�E�Ph�   �M��Q�l�����3҃} �U��}� uhD�j jh��j蓧������u̃}� u0�$����    j jh��ht�hD��q������   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U��E�Ph�   �M��Q�h���������t3�t	�E�   ��E�    �M܉M�}� uh̘j jh��j�x�������u̃}� u-�	���� "   j jh��ht�h̘�V������"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9�As
��A�E���M+M����U+щU؋E�Ph�   �M+M��U�D
P聦����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ����������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����������������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U��W�}3�������ك��E���8t3�����_��������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��������������������������������������̋�U��j������]���������������̋�U����E�    �E�    �	�E����E��}�$}Z�M��<�$MuK�U�k��°j�E��� M�M����M�h�  �U��� MP�D���u�M��� M    3��뗸   ��]��������������������������������������̋�U����E�    �	�E����E��}�$}O�M��<� M t@�U��<�$Mt3�E��� M�M��U�R�P�j�E�P�D������M��� M    ��E�    �	�U����U��}�$}3�E��<� M t$�M��<�$Mu�U��� M�E�M�Q�P�뾋�]��������������������������������������������������̋�U��j�hp/h�d�    P���SVW��A1E�3�P�E�d�    �E�   �=<_ u����j�A�����h�   �������E�<� M t
�   �   h  ht�jj�������E�}� u�I����    3��   j
�ڠ�����E�    �M�<� M uDh�  �U�R�D���u"j�E�P�ή����������    �E�    ��M�U�� M�j�E�P蝮�����E������   �j
������ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��E�<� M u�MQ�Y�������u
j蠳�����U�� MP���]�����������������̋�U��E�� MQ���]��������̋�U��EPj ���h�   �K�����]����������������̋�U��j�h�/h�d�    P�ĘSVW��A1E�3�P�E�d�    �} u3��   j莙������u3��oj�������E�    �EP�MQ�`l�е���URj �EP�MQ�UR�M�蛶���M��G����E�`l肫���E������   �j������ËE�M�d�    Y_^[��]��������������������������������������������������������������̋�U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� �����������������̋�U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]�������������������̋�U��j�h�/h�d�    P�ĘSVW��A1E�3�P�E�d�    �} u3��   j�Η������u3��pj�/������E�    �EP�MQ�`l�����U R�EP�MQ�UR�EP�M��ڴ���M�膵���E�`l������E������   �j�V�����ËE�M�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�M��M��v����M���,�k����E��l��l��l�} t�U��l�E��l���l    ��l    �M���,�xl�U��tl�E��l�M��l��l �E���]� ��������������������������������������������̋�U���H�M��M������M������=�l ��   ��l���?uG��l�B��@u8��l����l�U�R�ݠ����Ph���E�P�0�����P�M��s����v��l���?uS��l�H��$uEj �U�R� �����P�M��>����M��Q�����u��l��l�M�Q�j�����P�M�������U�R�S�����P�M�������M�������u	3��  �?�M��������t�֬����u��l���t��lR�M��h�����E�P�M�覑���=�l u2�M�趱������ljh`l��lQ覦�����E��U���l�=�l ��   ��lP��lQ�M�跪����l�U�E�E�M����tY�E���� u0�U���U�E��  �M���M�U���� u�M���M�����U�E��
�U���U�E���E�띋M�U����l��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M�jPh�l�M�胩����l��]���������������̋�U���h�a�����tH��l%������lj �M�Q�h�������l��    ��l�E�P�M�����E�  �  ��l���?�t  ��l����l��l���?uK��l�H��?u=�U�R謝������l���t��l����l��E�P�M莣���E�9  �M�Q�?������M��)����E�M������E��M��2�����u�U�R�M�L����E��  ��l�����   ��l���@��   �M�Q�Ƒ�����M���������   ��l��tn��l �E�P�M�Q�M��ٔ��P�M�聎����l���@t>�M�Q�q�����P�M��^����U�R�E�Ph��M�Q�M��ƞ����荔��P�M��5����)�U�R�E�Ph��M�Q�M�蛞�����b���P�M��
����}� t�M��ޡ���}� t�M��x����M�豟����u�M�財����t�U�R�M�$����E��   �   ��l���t��l���@ut��l���t��l����l臨����t:�}� u4�M��i�����u(�M��y���P�M�Q�|������U�R�M觡���E�U��E�P�MQ�Y������E�>�j�M�;����E�-�+��l���tj�M�����E��j�M�����E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�졀l���?uJ��l�B��$uj�MQ�Ǧ�����E�;�$��l����lj j �EP��������E��j j�MQ�������E]�������������������������������̋�U���h��A3ŉE䡀l���0�M�x5�}�	/��l����l�E�P�MQ�xl�����E�;  �6  �M��A�����l���?ubj �M�Q������P�M��	�����l���l����l��@t)��l����l��l�����ك�Q�M��ȏ���  jh ���lR���  ����u�E� ���l����l�9jh���lQ�ί  ����u�E����l����l��E�    �}� ��   �E�P讌�����9�����twj�M�Q�M�薣���U�R轪����P��l���EЃ}� t�E�P�M�豙���:h��M�袙��h��M�Q�U�R�E�P�M�Q腡�������K���P�M��U����:h��M��f���h��U�R�E�P�M�Q�U�R�I�����������P�M������N�E��t.��l���@u �M��x���P�M��\�����l����l�j@h�l�M��]���P�M��5����M��t�xl�#�����u�U�R�xl荈���E�P�M�]����E�M�3��|�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �M��=����M��5����E�    �E�    ��l��������l����l���������������_�o  �������|!�$�`!��l����lj�M�ɞ���E�  �M�趒���M����   �U�R�Ň����Pj<�E�P�)�����P�M������M��ۣ���ȃ�>u
j �M�詇��j>�M�蟇���} t�U���l���u�U�R�M腛���E�  ��l����l��l�M�j j �U�R�Q�����P�M������Eܣ�l�M�诘����u*��l�Q���1u�E�Pj~�M�Q�l�����P�M�趆���M��y�����u�U�R�M��2����E�P�M�����E�v  �%  ��l�Q�����P�M������  �E�   ��l�Q���t�P�M��������  ��l��������l����l���������������_��  �������"�$��!��l����lj�M������E��  ��l�B��� �Q�M��p����F  ��l�B��� �Q�M荆���E�  �  ��l�B��� �Q�M��f����M�������U�R�M輙���E�F  ��  jh���E�P��������M��p����M�Q�M舙���E�  ��l�B����Q�M������E��  ��l�B����Q�M�螔��j j �U�R������P�M��ф���M�蔖����u�M�������tj�M�ś���E�  �E�P�MQ�M������E�{  �  �  ��l�B����Q�M�������l���uj�MQ�M�蒃���E�4  ��l���0�E�x�}�rj�M�=����E�  �M�����R�M��������l��������l����l�����������������0�����������>  ������$�p"j �E�P�E������M�Q�UR�E�P��t���Qj ��|���R�M�赈�����Љ�����ɉ���E�^  �  �E�P�M�Q�M�謉��j,��d���R��l���P贅�������k���P�M��Ɋ��j,��T���Q��\���R茅�������C���P�M�衊��j,��D���P��L���Q�d�����������P�M��y���j)��4���Rj ��<���P������������P�M��O���j'�MQ�M��ڇ���E�  �;�U�R�EP�M������E�w  �!��l����lj�M膙���E�T  ��  ��l�B����Q�M��������  ��l��� �����l����l�� ��������������� t������0t!�N��l����lj�M�����E��  j h<��M�Q芃�����M������U�R�M�����E�  j�M�Ę���E�  �0  ��l���������l����l��������������������A������������	��   ���������"�$��"��l�Q���h�P�M�����E�  ��l�Q���h�P�M��������l���?u5��,���P�>�����P�M��z�����l���@u��l����l���$���Q�ٌ����P�M��E���h8��M��9����U�R�M�����E��j�M蝗���E�n�j�M茗���E�]�j�M�{����E�L�}� t
�M��4����-�M�������u!�E�Ph\������Q�������P�M��#����U�R�M�q����E��]ÍI ���-�  v���)Gi��
��  	

� ���% G         �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��Y}����l���l����l��@u��l���l����l��_tj�M�?����E�   ��l����lj �U�R�V�����j �E�P�H�������l���t��l���@t��l����l�ա�l���u��l����lj�M輒���E���l����l�M�Q�M�����E��]��������������������������������������������������������������������̋�U����   �M��=����E� �M��9�������  ��l�����  ��l���@��  ��l��t��l��u�E�P�M�,����E�(  �M�荌����uE�M�Qh��U�R�]�����P�M��z���E���t�M�Qj[�U�R�3�����P�M��}z���E� ��l���?�  ��l����l��l���@�����@�����$��@�����@���%��  ��@������)�$��)��l�B��_ua��l�Q��?uR��l����l�M�Q�U�Rj j �E�P��x������� ���P�M���y����l���@u��l����l�@�M�Q�U�Rj'�E�P�M�Q�������Pj`�U�R�/��������~��������P�M��ky����   ��l����l�M�Q�U�Rj j�E�P蕌���������P�M��1y����   j@h�l�M��<����M�Qh<��U�R輐����P�M���x���xl��|����u�E�P�xl�_x���w��l����l�U�R��|���Pj]�M�Qj j�U�R����������}������~��P�M��x���E��*�E�P��l���Q��t���R�����������~��P�M��hx���.�E�P��\���Qj j��d���R蜋�������~��P�M��8x��������l���<�����<��� t��<���@tW�W�M��Չ����tj�M��}���;�U�R��D���Ph���L���Qj��T����������P������~��P�M��w����
j�M��|���U�R�M������E��]Ð(A(R'�(�( �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����l���uj�M�e����E�T�R��l���?u3��l����lj �U�R�o�����Pj-�EP軅�����E��j �MQ�K������E��]�������������������������������������̋�U���   V�E�    ��l���Qu�E�X���l����l��l���uj�M藌���E�S  �N  ��l���0��   ��l���9��   �}� tG��l� ��/��E��U���l����l�U�R�E�P�M��܎��P�M�Q�U�R輌�����E��4��l� ��/��E��U���l����l�U�R�E�P�M�蕎���E��M��M�U�R�M�����E�  �  �E�    �E�    ��l���@��   ��l���uj�M萋���E�L  �W��l���A|7��l���P*�E��U���jz���ȋ��l���A���M��u��j�M�7����E��   ��l����l�e�����l���l����l��@tj�M������E�   �M��tX�}� t&�U�R�E�P�M��p���P�M�Q�U�R�_������E���E�P�M�Q�M��J����E��U��UЋE�P�M�ۇ���E�V�T�}� t&�M�Q�U�R�M��'���P�E�P�M�Q�������E���U�R�E�P�M������E��M��M��U�R�M胇���E^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����l���u3���   ��   ��l���0|8��l���9*��l���/�M���l����l�E��   �   �E�    ��l���@tY��l���u3��k�7��l���A|$��l���P�U�����l��T
��U������2��l����l뚋�l���l����l��@t�����E���]����������������������������������������������������������������������̋�U����   ��l���?u��l�B��$tj�M�����E�  ��l����l�tl�U��xl�E̋|l�M���\���蚑���M�蒑���M�芑����\����tl�E��xl�MЉ|l�M��{���M��{���E� ��l���?u/��l����l�U�Rj��T���P�eo����P�M��Dp���jj��L���Q胃����P�M��&p���M�������t��l�U���up��D���P�6p����Pj<��<���Q�����P�M��uw���M��I����Ѓ�>u
j �M��p��j>�M��p���E��t��l���t��l����l�M��tl�Ủxl�E��|l�M�Q�M�σ���E��]�����������������������������������������������������������������������������������������������������������������̋�U���|��A3ŉE��E�   �M���y����l�M���v�����  ��l����  ��l���@��  �}� t	�E�    �
j,�M���n����l���0�U�x4�}�	.��l����l�M�Q�U�R�|l�!s��P�M���u���  ��l�E�M��Hy����l���Xu��l����lh���M���}���%  ��l���$u7��l�H��$t)��l����l�E�P������P�M���m����   ��l���?��   �E�P�p�����}����tkj�M�Q�M�������U�R�#�����P��l���Eă}� t�E�P�M��}���.h��M�Q�U�Rh|��E�P����������}��P�M��3m���.h��M�Q�U�Rh|��E�P�Ǆ�������}��P�M��m����M��x��P�M�Q�r����P�M���l����l+U��~�|l��p����u�E�P�|l�5l���M�Q�M��?t���������l �U�R�M�����E�M�3��n����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ��A3ŉE血l��M���l����l�E�������������R��  ���������9�$��9�EP��m�����E�  ��l���@u$��l����lh���M�8l���E�S  �3��D���Q�~y����P�URh@���L����
l�����bq���E�  �EP�Ny�����E�
  �M�Q�Zm�����U�R�Nm�����M��|������   �M���{����t{jd�E�P�M��#�����uj�M轁���E�  �M��M��U���-u�E��E��E�.��E�.�M�Q�URje��4���P�M�Q��<����Pk�����o�����p���E�]  �j�M�T����E�I  ��x���R�l�����!z����tSj��h���P��x����x�����h���Q蜊����P��l����d�����d��� t��d���R�M��j���E��  �E���Du5h��MQ��x���Rh|���,���P�R��������z���E�  �3h��MQ��x���RhX���$���P����������y���E�m  �h  j j ��\���Q�|���������R�k������\���P�M�~}���E�/  j{��T����#����M�������������H|3������J~�(�����R�2w����P��T����kp��j,��T����i���E���������������F������������wx�������$�:�����P��j����P��T����p��j,��T�����h�������Q��j����P��T�����o��j,��T����h��������R�j����P��T�����o��j}�EP��T����Lm���E�-�+��l����lj�M����E�j�M����E�M�3��ii����]Ë�U9�5�5v677b6Q88s9 ��8�8"9�8�8���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �M��-q��詆���E��M�n���E��}���  uj�M�
}���E�  �B�}���  u�EPj�MQ�_y�����E�  ��}���  u�UR�M�
z���E�j  �E�% �  �0  �M��� �  t�U���   3���   ���������M��� `  ��Ƀ����������� t�U���   �� �����E�%   �� ����� ��� t>�M��� �  t�U���   3���   ���������
ǅ����    ������ ��
  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ t|�M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� @  tM�Di����t/��l����t&�U�R�{q����Pj �E�P�ys����P�M���c����M�Q�Uq����P�M�������U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t�E�%   ��������M���   ������������ �-  �U��� �  t�E�%   3�=   ���������
ǅ����    ������ ��   �U�R�w����P��|���Pj{�M�Q�M�h�����&i��P�M��bj���U�R�2n������}����u1hؤ��l���P�M�Qj,��t���R�Er�������s��P�M��j��hԤ�M��}���E�P�-f�����g����tR�f����tI�[}����u@�M�Q��T���Rj ��\���P�M�Qj ��d���R��q�������Qg�����lh��P�M��b���  �M��m���M��m���M��
m���M��m���M���l���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ �"  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t[�M���   ��   uJ��L���R觃����P�M��	a����D���P菃����P�M���`����<���Q�w�����P�M���`���k�U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t'�E�%   =   u��4���Q�
�����P�M��l`����,���R������P�M��T`���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t8�U��� �  t�E�%   3�=   ���������
ǅ����   ������ u;�\i����t��$���R��s����P�M��m_��������P��s����P�M��|���d����tO��b����t,�M�Q�����R�����P��b�������oe��P�M��_��������Q��b����P�M��N|���������R�b����P�M��4|���M�p����uA�M��p����u)��y����u �EPj ������Q�Zn����P�M��8f����UR�M��^���E�    �M��i���}� tNj ������P��i����PhФ������Q�v����P�M���e���Py����t�U�R�M�r���E��  �bj h`lj�Qs���������������� t�������i���������
ǅ����    �������E��M�Q������R�^i����P�M���]���E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ ��  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M���   ��   uzj,������R�E�P������Qj,������R�E�P������Qj,������R�E�Ph��������Q�rt��������a������b������a������b������a��P�M��&d���   �U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� tB�E�%   =   u3j,������Q�U�Rh��������P��s�������?a��P�M��c���h���M��v��hؤ������Q�M��gl��P�M��qc��j)��x���R������P�Cw����Pj(������Q�`k��������`��P�M��7c���U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� ��   �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t:�M��� �  t�U���   3���   ���������
ǅ����   ������ u�M�Q�M��eb���l����t��p���R�i����P�M��Db�����h���P�i����P�M���w���9]����t�}� t�M�Q�M��{Z���U�R�M��oZ���  �EP�M���a���M��� �  u.�U��� |  �� h  u�E�P�MQ�Zq�����E��	  �1  �U��� �  u,�E�% |  = p  u�M�Q�UR�_�����E�	  ��  �E�% �  u]�M��� |  �� `  uLhԤ�UR��X���P��j����P��P���Qj{��`���R�M���^������_�����j���E�N	  �  �E�% �  u.�M��� |  �� |  u�U�R�EP��h�����E�	  �[  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ thx��M��/s���  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ th<��M��ur����   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tI�M��� �  t�U���   3���   ���������
ǅ����    ������ th ��M��q���0�M��� �  u%�U��� |  �� x  u�E�P�M�Vk���E�  �M��� �  t�U���   3���   ����|�����M��� `  ��Ƀ���|�����|��� t�U���   ��x�����E�%   ��x�����x��� ��   �M��� �  t�U���   3���   ����t����
ǅt���    ��t��� u:�M��� �  t�U���   3���   ����p����
ǅp���    ��p��� t#�M�QhФ��H���R�m����P�M���U����E�P��@���Q�i����P�M���U���U��� �  t�E�%   3�=   ����l�����U��� `  ��҃���l�����l��� �x  �Hv�����R  �E�% �  t�M���   3ҁ�   ��h�����E�% `  �������h�����h��� t[�M��� �  t�U���   3���   ����d����
ǅd���   ��d��� t!�M�Qh����8���R�l����P�M���T���E�% �  t�M���   ��   �s  �U��� �  t�E�%   3�=   ����`�����U��� `  ��҃���`�����`��� t�E�%   ��\�����M���   ��\�����\��� �$  �U��� �  t�E�%   3�=   ����X�����U��� `  ��҃���X�����X��� t�E�%   =   ��   �M��� �  t�U���   3���   ����T�����M��� `  ��Ƀ���T�����T��� t�U���   ��   tU�E�% �  t�M���   3ҁ�   ��P�����E�% `  �������P�����P��� t2�M���   ��   u!�U�Rh���0���P��j����P�M��(S���t�����  �M��� �  t�U���   3���   ����L�����M��� `  ��Ƀ���L�����L��� tl�U��� �  t�E�%�   3Ƀ�@����H�����U���   3���   ����H�����H��� t&�M�Qhܣ��(���R�+j����P�M��nR���Z  �E�% �  t�M���   3ҁ�   ��D�����E�% `  �������D�����D��� tp�M��� �  t�U����   3����   ����@�����M���   3ҁ�   ��@�����@��� t&�E�Pḥ�� ���Q�wi����P�M��Q���   �U��� �  t�E�%   3�=   ����<�����U��� `  ��҃���<�����<��� tb�E�% �  t�M����   ��Ƀ���8�����U���   ��҃���8�����8��� t!�E�Ph�������Q��h����P�M��Q���U��� �  t�E�%   3�=   ����4�����U��� `  ��҃���4�����4��� t�E�%   ��0�����M���   ��0�����0��� t*�k����u!�U�Rh�������P�6h����P�M��yP���M���   t!�U�Rh�������P�
h����P�M��MP���M�Q�M�d���E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���x�E�    ��l���_u�U��� @  �U���l����l��l���A�  ��l���Z�  ��l���A�E���l����l�U��� �  �U��E���t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M�U����U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U��E��E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E܋M܉M��;�U��� �  t�E�%?����E���M��������M؋U؉U���E���  �E��k  �E����Eԃ}���   �M��$��_�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M̋ỦUЋEЉE����E���  �E��  �  ��l���$��  �E� ��l����l��l��Uȃ}�R�]  �E���`�$��_�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  ��l�Q��Pu��l����l��l����l��l��Eă}�Q��   �M���t`�$�``��l����l��g���  ��l����l��l���0|C��l���95��l���l�D
ѣ�l�g���E��M���   �M��E��-  ��E���  �7��l����l�Ng���	  �E���  �E���  �E���  �E���  ��  �E���  ��l����l��  �E���l����l��l���0|��l���5~$��l���t	�E���  ��E���  �E��z  ��l���0�E��M��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��M���t�U���    �U���E�%�����E��M����M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  ��l����l��  ��l���0��  ��l���8��  ��l��U졀l����l�M�������M��U�U��E���0�E��}��?  �M��$��`�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C��l���9u��l����l�E���  ���l���t	�E���  ��E���  �E���]ÍI �X Y�X Y�X YsX�Z�YG[^YuY�Y�Y�Y�Z�\ 																																																																					��ZZ6Z�Z�Z ��8]�]j^�^__3_G_Y_�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j �H����P�M���>����l���tl��l��E��l����l�U�U�}�0t�}�2t�}�5t(�5h���M��X���&�E�P�kP����P�M��E���j�M�wT���E�(�
j�M��A��hܤ�M���W���M�Q�M�Q���E��]���������������������������������������������������̋�U���@�M�� H��j j�E�P�1P����P�M���<���M���D����uN��l���tA��l���@t4�U�R�E�Ph��M�Q�U�R�?�������M������B��P�M��z<����l���@u��l����l�b��l���tj�M��KA���J�M��N����tj�M��3A���2�U�R�E�Ph��M�Qj�M��'S�����L�����RB��P�M���;���U�R�M�HP���E��]��������������������������������������������������������������������������̋�U�����l����  ��l���A�E���l����l�}���   j�M��iR���@������   �U�����U��}���   �E���4g�$�gj��E����P�M���J���|j�E����P�M��J���gj�E����P�M��J���Rj�E����P�M��J���=j�{E����P�M��oJ���(j�fE����P�M��ZJ���j�QE����P�M��EJ���U�R�M��N���E� �j�M�Q���E��j�M�yQ���E��]ÍI Kf`fuf�f�f�f�f�f ��������������������������������������������������������������������������������������������̋�U�졀l���@u"��l����l�EP�M�M���E���MQ�UR�":�����E]�����������������������̋�U��� �EP�M��YM����l��U��}� t�}�?tq�}�Xt��   �E�Pj�MQ�L�����E��   ��l����l�M���J����th���M��9���E�   ��E�Ph��MQ�P�����E�w��l����l�E�Kj �M���C��P�E�P�M�Q�U�R�g9����P�M��8���E�P�MQ�!>�����E�$�U�R�M��L���E��E�P�MQ��=�����E��]�������������������������������������������������������������������������̋�U���<�M��C����l��Mȃ}�B��  �U���4l�$� l�MQj�UR�UK�����E�j  h���M��dG���M�sI����u
j �M���7���EP�M���K����l����l�E�@��U�R�M��JJ��P�E�P�MQ�5=�����E�   ��l�B��$t<��l�Q��u�EPj�MQ�J�����E��  �j�M�&N���E�  ��l����l��l��Mă}�T�o  �U����l�$�xl��l����l�UR�EP�yV�����E�Y  ��l����lj�UR�EP�:�����E�0  ��l����l�E�Kj �M��vA��P�U�R�EP�M�Q�7����P�UR�M�����E��   ��   h���M���E���M��G����u
j �M��a6���EP�M��_J����l����l�E���U�R�M���H��P�E�P�MQ�;�����E�z��l����lj�M��L���E�\�G��l����lh��M�6���E�;�&�MQj�UR�
I�����E�"j�M�L���E��EP�MQ�3L�����E��]Ë��ij�i�il ��k�j�j�j\k9k�k�k�k ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� ��l��M�}�XtD�}�Zt�`��l����l�9����t	�E�����E� ��E�P�M�)4���E��   ��l����lh���M�4���E��   �U�R�6�����M��;������   ��l��M�}� t�}�@t`�}�Zt�v�U�R�M�!G���E�   ��l����l�a8����t	�E����E���M�Q�U�R�M��
C��P�M��F���E�>��l����l�M�Q�M�F���E� j�M�iI���E���U�R�M�F���E��]��������������������������������������������������������������������������������������������̋�U���,�E�   �M���<���M���9�����  ��l���@��   ��l���Z��   �}� t	�E�    �
j,�M���1����l�����   ��l���0�M�x3�}�	-��l����l�E�P�M�Q�tl��5��P�M��8���k��l�U�M��(<��P�E�P�6������l+M��~�tl��4����u�U�R�tl�Z0���E�P�M��d8����l;M�u
j�M���5���j�M���4���������U�R�M��D���E��]����������������������������������������������������������������������������������������̋�U���(��l���tg��l���Zu'��l����l�M��;��P�M�UD���E�^�0j)�UR�E�P�`K����Ph0��M�Q�G��������4���E�,�*j)�URj�E�Ph0��M��0������.������4���E��]�������������������������������������������������������̋�U���x��l����k  ��l��E���l����l�E� �E������M��+:���U��U��E���C�E��}��   �M����v�$��vh ��M��>���?  h���M��>���-  h���M��p>���  h��M��^>���	  h��M��L>����  hܥ�M��:>��hԥ�M��I����  �E����E���  ��l��U��E�E���l����l�U��U��}�Y�8  �E���,w�$��v�E������(  h̥�M��=���  hĥ�M��=���  h���M��=����   h���M��=����   h���M��v=����   h���M��d=���   h���M��R=���   h|��M��@=���   ��l����l�E�P�9����P�M��c-���M��&?����t�M�Q�M�A���E�~  �R�UR�E�P�D����Pht��MQ��D�����E�R  ��l����lj�M��2���hh��M��<���Qh���M��<���B��l����l�M�Q�g8����P�M��,���M��>����t�U�R�M��@���E��  �}����   �E��E��M���C�M��}���   �U����w�$��w�M�Qh\��U�R�D����P�M��I,���e�E�PhP��M�Q��C����P�M��),���E�U�U��E���E�E��}�w/�M����w�$��w�E�Ph\��M�Q�C����P�M���+���M�=����u�URj �E�P�q;����P�M��O3���M�Q�M�	@���E��   ��   �M��6���UR�M���?���}��uF�M��b+���E�P�M�Q�U�R��=�����M��>����uhh��M���E���E�P�M�?���E�}�M�=����tA�M���t$hH��M���:���U���th<��M��E����E���th���M��:���M�Q�U�R�EP�=�����E���MQj�UR�X>�����E��]Àr�r�r�r�r�r�r�r�ts�t   










	�I Vt,thszs�s�s�sVsJs�s�s�sqt 	
��&uuFu�u �I mu�u     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8��B����t�C����u	�E�   ��E�    �EЉE��M��3����l��U̡�l����l�M̉Mȃ}�Y��   �U����z�$��z��l����lhI��M�(���E�   h@��M��>7���kh4��M��/7���\h,��M�� 7���Mh ��M��7���>h��M��7���/��A���E��U�R��G����Ph��E�P��>����P�M��'���M��(2���}� t�M�Q�M��'���U�R��*����P�M��.���E�P�M�<;���E��]Ë��y�y�y�y!zzzPz ���������������������������������������������������������������������������������������������������������������������������������̋�U��EP��8�����E]����������̋�U����M���0����l�����   ��l��E�M��0�M�}�wH�U��$��|hl��M��5���>hd��M��5���/�-h\��M���4���hܥ�M���4���j�M�F<���E�~��l��M��l����l�E�E�M��1�M�}�w/�U����|�$��|�M�Qh\��U�R�<����P�M���$���E�P�M�9���E��j�M��;���E��]��{�{||||$|$|�|�|    ��������������������������������������������������������������������������������������������̋�U����   ��l���u�URj�EP�7�����E�  ��l���6|��l���9~ ��l���_tj�M��:���E��  ��l���6�U���l����l�}�)u[��l���t2��l���=�M���l����l�}�|�}�~�E�������EPj�MQ��6�����E�M  ��}� |�}�~�E������}��uj�M�':���E�   �M��.���UR�M��O7���E����  �M�Qh��U�R�:����P�M���"����l���t5�U�R�E�P�M�Q�%����Pj �U�R�I2��������(��P�M��"����E�Pj�M�Q�6����P�M��o"����l���t1��l���@u��l����l�j�M�Q9���E�J  ��M�Qj�UR�5�����E�.  ��+����t�E�P�s6����P�M���!����M�Q�\6����P�M��3?���U���tS�%'����t5�E�P�M�Q�U�R�]/����Pj �E�P�[1��������'��P�M��!����M�Q�0/����P�M���>����&����t)�U�R��x���P�M�Q�%%�������'��P�M��W!�����p���R�%����P�M��>���M� 3����u.j)��`���P�M�Qj(��h���R��0�������9&��P�M��!��j h`lj�!6������\�����\��� t��\�����+����0����
ǅ0���    ��0����E��M�Q�U�R�1,����j)��D���P��T���Q�<����Pj(��L���R�00�������%��P�M��(���A*����t�E���t�M�Q�M���'���1����t��<���R�2/����P�M���'�����4���P�/����P�M��l=���}� t�M�Q�M��	 ���j�M�7���E��U�R�M�F4���E��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����l�����   ��l���6|��l���9~��l���_un�UR�M��p���M�C0����u$�M�70����u�M��2����u�EP�M���%���M�0����u�MQ�M���%���U�R�EP��=�����E�   �>j �MQ�UR�EP�M�Q�������U�3Ƀ�*��Q�U�R�EP��!�����E�m�kj�M���4���MQ�M��]8���M�/����u�UR�M��D%���M�s/����u"�M�g/����u
j �M������EP�M��%���M�Q�M��1���E��]��������������������������������������������������������������������������������������������������̋�U���4�M��(����l����l��l��UЀ}�At�}�BtN�}�C��   �   �} u%�E����&u	�E�4���E���E�M̉��l����l�  �} tj�M�3���E�}  �E� j>�M��H7����l����l�N  �U�4���l����l�3  ��l���t��l�H��uj�M�&3���E�  �} tj�M�3���E��   ��l���0����l�Q�DЉE��l����l�}�v/j,�M��6���U�3�PR�M��e5��P�M�Q�M���!��P�M����j>�U�R�M�� ��P�M��u����l���$u��l����l�j^�E�P�M��v ��P�M��@����l���t��l����l�
j�M��M���M��,=���M�Q�M�`/���E��M�&���E��]�����������������������������������������������������������������������������������������������������������������������������������������������������̋�U���$  �M��]%���E� ��l����  ��l���$u8�MQ�U�R�EP�M�Q�'�����M���+����u�U�R�M�R.���E�  ��l���l�3҃�A����+��+ʉM�M���$���M���$���E�   �E艅����������t������tw��������   �  ������tW�2����tN�M��6+����u/j�$����P�M�Qj �U�R�M��w������)��P�M��:���j��#����P�M���(���   �k����tN�M���*����u/j
�#����P�E�Pj �M�Q�M�������h)��P�M������j
�#����P�M��}(���`�����tN�M��*����u/j	�_#����P�U�Rj �E�P�M��������)��P�M�����j	�0#����P�M��$(����E�    �}� t|��l����l��l���$u8�MQ�U�R�EP�M�Q�'%�����M���)����u�U�R�M�n,���E�  ��l���l�3҃�A����+��+ʉM�}� �)�����l���t��l����l�}���  �EP�M�����M�Q�U�R�M�����P�M�����M��T)����u)�E�P��|���Qj �U�R�M���������P�M��\���M��)����u,�E�P��l���Qj ��t���R�M��a�����|��P�M��$���E���  �} tj�M�.���E�  �M���tz�E�Ph���d���Q�.����P�M�������l���t,�M�Q��T���R��\���P�����������P�M������M�Qj��L���R�*����P�M��~���$��l���t��D���R�k����P�M��3����l���uj�M��u���/��l���l����l��@tj�M�/-���E�  �\����t[�U��������������t�B�} tj�M��,���E�t  �E�P��4���Q��<���R�_#���������P�M�����#�E����u��,���Q�3#����P�M���2���U��t!�E�Ph|���$���Q�-����P�M��a���U��t!�E�Pht������Q��,����P�M��8���} ��   �M��&������   �M�)����u�M��&����t:�M�E(����t�UR�M�������EPj �����Q�$����P�M��b���@�UR������Pj �����Q�URj �����P�P$����������������P�M�� ���*�M�M&����u�MQj ������R�$����P�M������M��6'���E���t�M��)$���M�Q�M�(���E��   �j�M�>+���E�   �   �} ux�M��%����ul�M�(����u�M��%����t�URj�EP�o'�����E�u�9�MQ�URj ������P�MQj������R�B'�����������������E�:�8�} u%�M�Z%����u�EPj�MQ�	'�����E��j�M�~*���E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����l����  �} t]��l���XuO��l����l�M�%#����th���M�9���E��   ��URh��EP��(�����E��   ��l���Yu%��l����l�MQ�UR�v�����E�   �EP�M�Q�'�����M�����t �U�Rh���E�P�r(����P�M�����*�M��%����t�M�Qh���U�R�F(����P�M�����E�P�M��$���E���MQj�UR��#�����E��]��������������������������������������������������������������������������������̋�U���   ��l����s  �����E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M���(��������������P�MQ�&�����E�  �  �M�����M��"����thh��M��*���M�� ����tR�U��E����E���tB��l���t5j]�E�Pj �M�Q�$����Pj[�U�R���������R��P�M����뢋M�� ����u^�M�M"����t�E�P�M�Q�M�A��P�M������7�U�R�E�Pj)�M�Q�URj(�E�P�t���������������P�M�����M�Q�U�R�>�����M��z���E�P�M��"���E�   �   �M�B ����uSj]��|���Qj�U�Rh���E�P�MQj(�U�R���������������}�����a��P�EP�%�����E�?�=j]��d���Qj��l���Rj[��t����'�����<����� ��P�EP��$�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j'�EPj �M�Q�"����Pj`�U�R���������H���E��]�����������������������̋�U����E��Kj�M�����P�E�P�M�����P�MQ������E��]����������������������̋�U��Q�E�T��E�P�MQ�UR�EP� �����E��]��������������������̋�U��Q�E��K�E�P�MQ�UR�EP�s �����E��]��������������������̋�U��EP�MQ�UR�EP�; �����E]��������������̋�U��j�EP�<!�����E]��������̋�U��j �EP�!�����E]��������̋�U��j �EP�� �����E]��������̋�U��EP�MQ�"�����E]������̋�U��Q��l��M��}� t)�}�At�0��l����lh���M�3���E�j�M�J"���E�j�M�;"���E��]���������������������������������̋�U���@�EP�M��C���M�������b  ��l����Q  �E�P�M�Qj �U�R�E�P�p����������������P�M��
���M�������  ��l���@��   h���M���$���M��������   ��l�����   ��l���@txj'�M�Q�U�R�2����Pj`�E�P���������?��P�M������l���@u��l����l�M������t��l���@th���M��\$���Z����M�������t ��l���u
j�M�����j}�M���	����l���@u��l����l�'�M������t�U�Rj�E�P������P�M��P	���M�Q�M����E��]����������������������������������������������������������������������������������������������������������������̋�U��EP��	�����E]����������̋�U����E��Kj �M����P�E�P�M����P�MQ�E	�����E��]����������������������̋�U����EP�M����h���M���"���M�Q�:����P�M����j}�M��m����l���@u��l����l�U�R�M�N���E��]��������������������������������̋�U���,j h`lj�������E��}� t�M�����E���E�    �EԉE�M�Q�U�R������EP�M�Qj �U�R�E�P�)��������������P�M��P���M�Q�M����E��]������������������������������������������������̋�U�졐l�������]����������̋�U�졐l%   �����]��������̋�U�졐l�������]����������̋�U�졐l�������]����������̋�U�졐l�������]����������̋�U�졐l��`3Ƀ�`����]�������̋�U�졐l%�   �����]��������̋�U�졐l%   �����]��������̋�U�졐l%   �����]��������̋�U�졐l%   ]���������������̋�U�졐l%    ]���������������̋�U�졐l% @  ]���������������̋�U�졐l% �  �����]��������̋�U�졐l%   �����]��������̋�U�������t�E��(����M��(���]���������������������̋�U�졐l�������]����������̋�U��EP�MQ�`l����]�������̋�U����M�E������E�} t�MQ�U��Ѓ���   ��   �} w�E   �M�Q;U��   �}   v3��   jh`lh  ������E��}� t�M��!���E���E�    �E��E��}� tA�M�y t�U�B�M���U�E��B��M�U��Q�E�M��H�   +U�E�P�3��!��M�Q+U�E�P�M�Q�E�H�D
��]� ���������������������������������������������������������������������̋�U��Q�M��E��     �E���]�������̋�U����EP�MQ�UR�M��T�����	���E��]���������������������̋�U����EP�MQ�UR�M�������I	���E��]����������������������̋�U����EP�MQ�UR�M�������		���E��]����������������������̋�U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]�����������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M������E���]� ������������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��} tdj h`lj�z�����E��}� t�EP�M������E���E�    �M��U��E����Ƀ�������   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ���������������������������������������������������������������������������������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ��"  ���E��}� v�U�R�EP�M������E���]� ���������������������������������������������������������������������̋�U���V�M�E�H�� ����U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E��     �M�Q�������E�P�M�Q�������E�P�M�Q�������E�P�M�Q������E�P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	������t�U����U���E�H�� ������U�J�   ������E�P�M�Q�M�����U����t<�U�E���M�	���u�;�t�U�B% ������M�A�U��    �!�M��q����u�E�H�� ������U�J��E�H�� ������U�J��E�H�� ������U�J�E�^��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�졐l%   ]���������������̋�U���$��A3ŉE��M܍E��E��M܋Q�� ����E܉P�M��    �U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%����M܉A�U�� �E����E�j j
�MQ�UR�����0�� �M��j j
�UR�EP����E�U�MMu��U��E�+й   +�Q�U�R�M������E܋M�3�������]� ����������������������������������������������������������������������������������������̋�U���(��A3ŉE��M؍E��E܋M؋Q�� ����E؉P�M��    �U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%����M؉A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U܃��U�j j
�EP�MQ������0�� �U܈j j
�EP�MQ�d���E�U�UUu��E��t�M܃��M܋U��-�E܍M�+��   +�R�E�P�M�����E؋M�3�������]� ��������������������������������������������������������������������������������������������������������̋�U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�������M���U��: u�E��H�� ������U��J�E���]� �����������������������������������������������������������������������̋�U��Q�M��E��H����3�������]���������������̋�U��Q�M��E�3Ƀ8 ������]������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J�E���]��������������̋�U��Q�M��E��@������]�������̋�U����M��M��U����u�E��H��	��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��M������u�E��H��   �U��J��]���������������������̋�U����M��M�������u�E��H��
��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��    �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� @  �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� �  �U��J��]�����������������̋�U��Q�M��M�������t3���E���U����ȋ�Ћ�]�����������������̋�U��Q�M��M������t2���E���U����ȋB�Ћ�]����������������̋�U����M�M��e����uX�} u*�M�������Ej h`l�EP������E��M��M�} t �U�E�L�Q�UR�M������E��E��  ��} t�M� �E��]� �������������������������������������������̋�U��Q�M��M������t�E��EP�MQ�U���M��	��B�Ћ�]� ����������������������̋�U����M�E�P�M������MQ�M�������U�R�M�����E��]� ����������������������̋�U����M�E�P�M�����MQ�M���
���U�R�M����E��]� �����������������������̋�U����M�E�P�M��P���MQ�M��~����U�R�M�8���E��]� �����������������������̋�U����M�E�P�M�� ���MQ�M������U�R�M�����E��]� �����������������������̋�U����M�E�P�M�����MQ�M��}����U�R�M����E��]� �����������������������̋�U����M��} t_j h`lj�*�����E��}� t�EP�M��R�M��6���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ������������������������������������̋�U����M��M�������tb�E��tZ�M�� ����t�MQ�M��	���?j h`lj�Q�����E��}� t�UR�M��	���E���E�    �E�P�M������E���]� ���������������������������������������������̋�U����M��M��������tu�} to�E���te�M��Y�����t�UR�M��2����Kj h`lj������E��}� t�EP�  ��P�MQ�M��a����E���E�    �U�R�M��	���E���]� ������������������������������������������̋�U��Q�M��M�������tG�M������t�M�����P�M�������(�M�������t�EP�M�������M�R�M��y���E���]� ��������������������������̋�U����M��M���������   �} ��   �M�������t�EP�M��!����j�M�Q�����t�M�E�����u@j h`lj�C�����E��}� t�MQ�M������E���E�    �U�R�M������M�����P�M������E���]� ���������������������������������������������̋�U��Q�M��M�������tC�M��K�����u�}t�}u�EP�M��i�����} u��MQ�A
����P�M�����E���]� ������������������������������̋�U����M��M��%�����t3�M�-�����u'�M�����E��E�%�   �M��Q�� ���ЋE��P�E���]� ���������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M�������E���]� ������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�  ��P�UR�M������E���]� ���������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h`lj�������E��}� t�MQ�M������E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������̋�U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ�	�����U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ������������������������������������������������������������������̋�U����M�E�8 tj�M������  �} ��   �} ��   �M�M��}� t�}�t�u�U�B% ������M�A�   j h`lj�X������E��}� t�U�P�M�� ���E���E�    �M�U��E�8 u�M�Q�� ������E�P�[j h`lj��������E��}� t�MQ�UR�M�������E���E�    �E�M��U�: u�E�H�� ������U�J��E�H�� ������U�J��]� ����������������������������������������������������������������������������������������̋�U��Q�M��E�3Ƀ8	������]������̋�U��Q�M��E�� �����E���]�������̋�U����M�M�������uf�M�y�����uZj h`lj��������E��}� t�EP�M�������E���E�    �M��M��}� t�U����M��U��M�U��T��E��]� �����������������������������������������̋�U��Q�M��} |�}	~j�M�����E�;�9�E��8�t
�M��U;~j�M������E���E�M��T�R�M�����E��]� ��������������������������̋�U��Q�M��E�� ���E���]�������̋�U��Q�M��M������E�� Ц�M��U�Q�E���]� �������������������̋�U��Q�M��   ��]��������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E;Es�M�U��B��M���M�E��]� �����������������̋�U����M��M�������E�� ��} tP�} tJj h`l�MQ�������E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ�S  ����U��B    �E��@    �E���]� ������������������������������������������������̋�U��Q�M��E��@��]�������������̋�U����M��E��x t�M��Q�E��H�T
��U���E� �E���]����������������������������̋�U��Q�M��E��HQ�U��BP�MQ�UR�[������]� ������������������̋�U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�"  ���EE��]���������������������̋�U����M��M��<����E�� ��} t#�M�������t�M�������u	�E�    ��M�M��U��E��B�E���]� ����������������������������������̋�U����M��E��x t�M��I�����E���E�    �E���]��������������̋�U����M��E��x t�M��I�����E���E� �E���]�����������������̋�U����M��E��x t�MQ�UR�E��H�a����E���M�M��E���]� ��������������������̋�U��Q�M��M�������E��  ��M��U�Q�E��H����Ƀ�����U��J�E���]� ��������������������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E��x��,"���]�����������������̋�U��Q�M��E��xujh��MQ�UR���������E��]� ���������������������������̋�U��j�hn�
d�    P��A3�P�E�d�    �Dm��uM�Dm���Dm�E�    j �m�H���j�m�<���j� m�0���j�,m�$����E������} |�}}�Ek�m��,m�M�d�    Y��]��������������������������������������������������������̋�U��Q�M��M������E�� ��M��U�Q�E��M�H�U��B�����E���]� ����������������̋�U��QV�M��E��x }.�M��Q�E��H���Ћ��M��Q�E��H������M��q�U��B^��]��������������������̋�U����M��E��H�U��B��ȋB�ЈE��M���u�U��B�M��I��B�ЈE��E���]������������������������̋�U����M��EP�MQ�U��B�M��I��B�ЉE��M�;Ms�UR�E�P�M��Q�E��H��B�����E���]� ����������������������̋�U��Q�E�    �	�E���E�M���t�E����E���E���]����������������������������̋�U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]��������������������������̋�U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]������������������������̋�U��Q�E�    �}�wC�EP�9������E��}� t�*�=@_ u�*����    ��MQ�u�������u����UR�_�����������    3���}� u������    �E���]���������������������������������������̋�U��Q�=<_ u�����j�D�����h�   �������} t�E�E���E�   �M�Qj �<_R�����]�������������������������̋�U��QV�E�    �} u�4�EPj �<_Q����E��}� u�$�P�Q�������������0^��]����������������������������������SVW�T$�D$�L$URPQQhP�d�5    ��A3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�����   �C�����d�    ��_^[ËL$�A   �   t3�D$�H3�����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�����3�3�3�3�3���U��SVWj Rh��Q����_^[]�U�l$RQ�t$������]� ���������������������������������������������������������������������������������������������̋�U��E�Hm]�����������������̋�U��Qj�������HmP�ܑ�E��MQ���Hmj��������E���]�����������������̋�U��} th��j jWh(�j���������u�j �3�����]���������������������������̋�U��HmP�ܑ]�������������̋�U��Q�HmP�ܑ�E��}� t�MQ�U�����u3���   ��]��������������������������̋�U��   ]����̋�U���0�    ]���������������̋�U���V3��} ���E�}� uhT�j jHh�j���������u̃}� u-�~����    j jHh�h��hT��������3��   �}�v�K����    3��~�} u�E   �URj �<_P�̒�E��MQ�URj�<_P�Ȓ�E��}� u:�}� @  w�M;M�w�x   ��t�U�U���$�P��������������0�E�^��]����������������������������������������������������������������������������̋�U����E�����j j�E�Pj �<_Q�В��t�}�u	�E�   ��E�    �E���]�������������������������̋�U���V�E�E��} u�MQ���������   �} u�UR�f�����3��   �E�    �}�w)�} u�E   �EP�MQj �<_R�Ȓ�E���EP������������    3��e�}� u	�=@_ u%�}� t��$�P���������U����0�E��1�MQ��������u�$�P���������(����03���J���^��]����������������������������������������������������������������������̋�U��Q�E�����j j �<_P�0���u�E������E���]�����������������̋�U���^���]����̋�U���<�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� uhoj jih��j��������u̃}� u.�����    j jih��h��ho�h���������  3Ƀ} ���M̃}� uhx�j jnh��j�&�������u̃}� u.�����    j jnh��h��hx�����������   �E�E��M��A����U��BB   �E�M�H�U�E��M�Qj �UR�E�P�k������E��} u�E��Q�M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj �������EċE���]��������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�=�������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ���������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��������]��������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�T�������]������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP��������]����������������̋�U��Q�E�E��M�Qj �UR�EP�MQ���������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��������]��������������������̋�U��Q�E�E��M�Q�UR���������]����������������̋�U��Q�E�E��M�Q�UR�M�������]����������������̋�U��Q�E�E��M�Q�UR�EP� �������]������������̋�U��Q�E�E��M�Q�UR�EP���������]������������̋�U��E��=   vh��j j8h0�j�6�������u̋UR�EPj �9�����]����������������������������̋�U����EP�M�������M����   vh��j jDh0�j���������u̃}�|5�}�   ,�M������ ���   �U�Q#E�E�M�������E��1�'�M����������   �B�#E�E�M������E���M�������]��������������������������������������������������̋�U���(�EP�M�������}�|6�}�   -�M��W�������   �E�B#M�M��M��.����E��   �M��*���P�U�����   R�)�������t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M������� �HQ�M��������BP�M�Q�U�R�E�Pj�M�����P������ ��u�E�    �M������E���M�#M�M؍M��k����E؋�]������������������������������������������������������������������������������̋�U��=�m u�E�K�A#E��j �UR�EP�,�����]���������������������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�,�����   u������r)��$����Ǻ   ��r����$���$� ���$�����@�d�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$����� ���(��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�<��I �Ǻ   ��r��+��$����$�����������F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I @�H�P�X�`�h�p����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]���������������������������������̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�������������������������������������������̋�U��j�h 0h�d�    P���SVW��A1E�3�P�E�d�    �e��E�   �E�    �E�P��������u�E�    �E������E��   �M+M�M܋U�R�E�P�������E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]������������������������������������������������������������������������������̋�U��h�����Lm]���������̋�U��j�h 0h�d�    P���SVW��A1E�3�P�E�d�    �e��w����@x�E�}� t#�E�    �U��E�������   Ëe��E�����������M�d�    Y_^[��]��������������������������������̋�U��Q�����@|�E��}� t�U��q�����]�������������̋�U��j�h@0h�d�    P���SVW��A1E�3�P�E�d�    �e�LmP�ܑ�E�}� t#�E�    �U��E�������   Ëe��E�����������M�d�    Y_^[��]��������������������������������������������̋�U��E�Pm�M�Tm�U�Xm�E�\m]�����������������������̋�U��j�h`0h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    �}t�}u�T  �}t�}t�}t�}t
�}�F  j �������E�    �}t�}u=�=`m u4jh���Ԓ��u�`m   ��$���� ����0�E�   �E�E̋M̃��M̃}���   �U������$�|��PmQ�ܑ�E�}t�UR���Pm�r�TmP�ܑ�E�}t�MQ���Tm�L�XmR�ܑ�E�}t�EP���Xm�%�\mQ�ܑ�E�}t�UR���\m�E������   �j �������Ã}� t��   ��   �}t�}t�}t��   �9����E؃}� u��   �E؁x\`muLhY  h��j��mQ�������EȋU؋EȉB\�}� t��mQh`m�U؋B\P���������j�M؋Q\R�EP�5  ���E��}� u�L�M��Q�U�}t5�E��H;Mu*�U��E�B�M����M���mk��E�P\9U�r��ˋE��   �M�MċUă��Uă}�w�E������$�������x3�t	�E�   ��E�    �E��EЃ}� u!hl�j h�  h��j���������u̃}� u.�V����    j h�  h��h�hl���������������M�d�    Y_^[��]Ë��d���>��� �I ����     ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h�0h�d�    P���SVW��A1E�3�P�E�d�    j �N������E�    �} u�E�Pm�E܋Q�ܑ�E��E�   ��E�Tm�U܋P�ܑ�E��E�   �}� t�}�t
�-����M܉�E������   �j �`�����Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������̋�U��j�h�0h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U������$����E�Pm�MЋ�U�E؃��E��  �E�Tm�MЋ�U�E؃��E���   �E�Xm�MЋ�U�E؃��E���   �E�\m�MЋ�U�E؃��E��   �{����E��}� u�����  �M��Q\R�EP��  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!hl�j h�  h��j���������u̃}� u1�Z����    j h�  h��h��hl�����������4  �E�P�ܑ�E�}�u3��  �}� uj�<����}� t
j �������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<��m�M��	�Uԃ��Uԡ�m�m9E�}�M�k��U��B\�D    ���
�L����MЉ�E������   ��}� t
j �y�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë�:���t���W��� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��Q;Ut�E����E���mk�M9M�s�ً�mk�U9U�s�E��H;Mu�E���3���]������������������������������������̋�U��XmP�ܑ]�������������̋�U���������d]�����������������̋�U��������`]�����������������̋�U��E�hm]�����������������̋�U���$V�hmP�ܑ�E�3Ƀ} ���M��}� uh�j jDh��j��������u̃}� u0�����    j jDh��h��h���������   �  �E�     �}� �_  h|�� ��E�}� ut3�t	�E�   ��E�    �U��U�}� uh �j jPh��j�s�������u̃}� u0�����    j jPh��h��h ��Q������   ��   h��M�Q����E��}� ��   3�t	�E�   ��E�    �E܉E�}� uh �j jVh��j��������u̃}� uD�$�P���������c����0j jVh��h��h ��������$�P�������V�U�R���E������E��E�Phhm�ؒ;E�t
�M�Q���j�UR�U���u������    ������ �3�^��]����������������������������������������������������������������������������������������������������������������������������������������̋�U��jj �EP�MQ��  ��]���������������������̋�U��jj �EPj ��  ��]�������̋�U��jj �EP�MQ�  ��]���������������������̋�U��jj �EPj �|  ��]�������̋�U��jj �EP�MQ�Z  ��]���������������������̋�U��jj �EPj �,  ��]�������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj ��  ��]��������������������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj �y  ��]��������������������̋�U��jh  �EP�MQ�G  ��]������������������̋�U��jh  �EPj �  ��]��������������������̋�U��jhW  �EP�MQ��  ��]������������������̋�U��jhW  �EPj �  ��]��������������������̋�U��jj�EP�MQ�  ��]���������������������̋�U��jj�EPj �\  ��]�������̋�U��jj �EP�MQ�:  ��]���������������������̋�U��jj �EPj �  ��]�������̋�U��jj �EP�MQ��   ��]���������������������̋�U��jj �EPj �   ��]�������̋�U����EP�M������M�薸���x t8�M�舸���H�y�  u$jj �UR�EP�i   ���E�M��Q����E���E�    �M��=����E��]��������������������������������̋�U��j �EP蚷����]�����������̋�U��j�h��
d�    P����A3�P�E�d�    �EP�M��P����E�    �M�M�M�蹷���P�E�L#Mu;�} t�M�蛷������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M��F����E��M�d�    Y��]��������������������������������������������������������������̋�U����} uh`�j jdh�j�z�������u̋M�M��U�R�q������E��E��H��   u$������ 	   �U��B�� �M��A����G  �-�U��B��@t"����� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6������� 9E�t�������@9E�u�M�Q��������u�U�R�{������E��H��  ��   �U��E��
+Hy!hP�j h�   h�j���������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�:������E��q�}��t!�}��t�M����U���������U���E�B�E��H�� t7jj j �U�R�1������E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P蜴�����E�M�;M�t�U��B�� �M��A�����E%�   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   ��A3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M�达���E�    �q����E�3Ƀ} �������������� u!h��j h  h�j虳������u̃����� uF�'����    j h  h�h��h���q�����ǅ ��������M������� �����  �E�������������Q��@��   ������P�)������������������t-�������t$���������������������������
ǅ���B������H$�����х�uV�������t-�������t$���������������������������
ǅ���B������B$�� ���ȅ�tǅ ���    �
ǅ ���   �� ��������������� u!h��j h  h�j�$�������u̃����� uF�����    j h  h�h��h���������ǅ��������M��0���������U  3Ƀ} �������������� u!hoj h  h�j蜱������u̃����� uF�*����    j h  h�h��ho�t�����ǅ��������M������������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���g  ������ �Z  �������� |%��������x��������x����������
ǅ����    ���������������������������������������������������������  �������$���E�    �M�路��P������R軱��������   ������P�MQ������R�t  ���E��������U���U����������؉�����u!h��j h�  h�j�ݯ������u̃����� uF�k����    j h�  h�h��h��������ǅ��������M������������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK����������$���E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�	������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�������Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ����������$���E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ��������P�$��U���0  u�E�   �E��M���  tUǅ|���    �UR诽����f������������Ph   ������Q�U�R�$�������|�����|��� t�E�   �&�EP������f��x�����x����������E�   �������U��W  �EP�W�������t�����t��� t��t����y u��N�U��E�P�;������E��P�M���   t&��t����B�E���t�����+����E��E�   ��E�    ��t����B�E���t�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������l����MQ�������E��U���  te�}� u��N�E��E�   �M���h�����l�����l�������l�����t��h������t��h�������h����ɋ�h���+M����M��[�}� u	��N�U��E���p�����l�����l�������l�����t��p������t��p�������p����ɋ�p���+E��E��  �MQ��������d���蒷������   3�tǅ����   �
ǅ����    ��������`�����`��� u!h@�j h�  h�j��������u̃�`��� uF�u����    j h�  h�h��h@�迼����ǅ��������M������������  ��  �U��� t��d���f������f����d�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h�j�Ú�]  R�������E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���X�����\����M�����P�E�P�M�Q������R�E�P�M�Q��X���R��AP�ܑ�Ѓ��M���   t$�}� u�M�薧��P�U�R��AP�ܑ�Ѓ���������gu*�U���   u�M��a���P�E�P��AQ�ܑ�Ѓ��U����-u�M���   �M��U����U��E�P�1������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�M�������H�����L����   �U���   t�EP�%�������H�����L����   �M��� tB�U���@t�EP�)���������H�����L�����MQ�����������H�����L����=�U���@t�EP���������H�����L�����MQ�̽����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��M̋Ũ��U̅���@����D���t{�E��RP��D���Q��@���R�6�����0��T����E��RP��D���P��@���Q蘽����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �J  ���U�R������P�MQ�U�R�E�P�{  ���M���t$�U���u������P�MQ��<���Rj0��  ���}� ��   �}� ��   ǅ$���    �E���8����M܉�4�����4�����4�������4�������   ��8���f�f������������Pj��(���Q��0���R�5�������$�����8�������8�����$��� u	��0��� uǅ���������*�M�Q������R�EP��0���Q��(���R�z  ���V�����E�P������Q�UR�E�P�M�Q�T  �������� |$�U���t������P�MQ��<���Rj ��  ���}� tj�E�P�������E�    �v���������������M��ּ��������M�3��s�����]Ì�����0�}������
������"�+� �I 8���	���� ���D���^����Z�<���W��NjE   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP蝯�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A�]��������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��E����U�
�E�f�A�]�������������������̋�U����E�    �E�E�}� |,�}�~�}�t��T]�M��U�T]�y�T]�E��o3�t	�E�   ��E�    �U��U��}� uhP�j j9hذj衙������u̃}� u+�2����    j j9hذh��hP������������E���]���������������������������������������������������̋�U��E�X]]�����������������̋�U���@��A3ŉE��E�    �u����E��E�    �E�    �E�    �=lm ��   h�� ��Eԃ}� u3��  h���E�P����E��}� u3��  �M�Q���lmh��U�R���P���pmẖ�E�P���P���tmh���M�Q����E��U�R���|m�=|m th���E�P���P���xm�xm;M�th�|m;U�t]�xmP�ܑ�EЋ|mQ�ܑ�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�pm;M�t�pmR�ܑ�Eȃ}� t�UȉE�}� t*�tm;E�t �tmQ�ܑ�Eă}� t
�U�R�UĉE�lmP�ܑ�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��������]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uhh�j jh�j��������u̃}� u0詯���    j jh�hвhh���������   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E��M���Qh�   �U��R�(�����3��} ���E��}� uhD�j jh�j�O�������u̃}� u0�����    j jh�hвhD��-������   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E܋M���Qh�   �U��R�/����������t3�t	�E�   ��E�    �U؉U�}� uh(�j j h�j�?�������u̃}� u0�Э���    j j h�hвh(��������   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���MԋU���Rh�   �E��P����������t3�t	�E�   ��E�    �EЉE�}� uh̘j j*h�j�+�������u̃}� u-輬��� "   j j*h�hвh̘�	������"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�As��A�U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�1�����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uhh�j jh�j��������u̃}� u0谪���    j jh�h̳hh���������   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E�M���Qh�   �U��R�3�����3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���M��U���Rh�   �E��P�ʐ����3Ƀ} ���M��}� uhD�j jh�j��������u̃}� u0肩���    j jh�h̳hD��Ϣ�����   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}������t&�M;Mrh�j j+h�j�C�������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E܋M���Qh�   �U��R����������t3�t	�E�   ��E�    �U؉U�}� uh̘j j>h�j�.�������u̃}� u-迧��� "   j j>h�h̳h̘�������"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9�As��A�M���U+U����E+EԋM���Qh�   �U+U��E�LPQ�4�����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���E����E���t��E�+E������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uhh�j jh��j��������u̃}� u0�y����    j jh��hh�hh��ƞ�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E�M���Qh�   �U��R�������3��} ���E��}� uhD�j jh��j��������u̃}� u0谤���    j jh��hh�hD���������   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���M��U���Rh�   �E��P����������t3�t	�E�   ��E�    �E܉E�}� uh̘j jh��j���������u̃}� u-萣��� "   j jh��hh�h̘�ݜ�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9�As��A�U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR������3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�j jh�j�/�������u̃}� u0������    j jh�h��h��������   �J  �} u\�U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U�E�Ph�   �M��Q�G�����3���  �} ��   �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U��E�Ph�   �M��Q������3҃} �U��}� uhD�j jh�j��������u̃}� u0虠���    j jh�h��hD��������   �#  �M�M��U�U��}�u5�E��M���E���U����U��E���E��t�M����M�t���y������t&�U;Urh�j j+h�j�\�������u̋M��U���M���E����E��M���M��t�U����U�t�E���Et�} u�M�� �}� ��   �}�u�UU�B� �P   �?  �E�  �}�tI�}���t@�}v:�M��9�As��A�U��	�E���E܋M�Qh�   �U��R�B���������t3�t	�E�   ��E�    �U؉U�}� uh̘j j>h�j�R�������u̃}� u-����� "   j j>h�h��h̘�0������"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9�As��A�M���U+U����E+EԋM�Qh�   �U+U��E�LQ�Z�����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M��o����MQ�UR�EP�MQ�M��ւ��P�.   ���E�M�趝���E��]�������������������������̋�U����E�    �E��Q�U�j j �EP�MQ����E�}� u3���   �}� ~63�u2�����3��u��r#h��  �E�L Q�P�����P�������E���E�    �U�U��}� u3��s�E�P�M�Q�UR�EP�����u�H�F�} uj j j j j��M�Qj �U�R���E��!j j �EP�MQj��U�Rj �E�P���E��M�Q�~������E���]��������������������������������������������������������������������������̋�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�f������.�}���  t%3�u!h�j h�   h��j�d�������u̋�]��������������������������̋�U���$�} t�} v	�E�   ��E�    �E�E��}� uhh�j jh��j���������u̃}� u0艚���    j jh��ht�hh��֓�����   �(  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9�As��A�U��	�E+E��E�M���Qh�   �U��E�PQ�"����3���   3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E��M���Qh�   �U��R��~��������t3�t	�E�   ��E�    �U܉U�}� uh̘j jlh��j��}������u̃}� u-�c���� "   j jlh��ht�h̘谐�����"   ��   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E�}� v�M����t�E���E�M���M��܋U����:u2�} t!�}s�  j�MQ�UR�EP�˒�����M���M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E؋M���Qh�   �U��R��{�����E�    �E�    �E�E��	�M���M�U����t4�M����/t�E����\u�U���U���E����.u�U�U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR�ȑ�����E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9�As��A�M��	�U���UԋE���Ph�   �M��Q��z�����}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR�������}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R�������   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR謐�����}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9�As
��A�E��	�M(���MЋU���Rh�   �E$��P��y����3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9�As��A�M��	�U���ŰE���Ph�   �M��Q�Vy�����} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���EȋM���Qh�   �U��R��x�����} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9�As
��A�E��	�M ���MċU���Rh�   �E��P�x�����}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9�As��A�M��	�U(���U��E���Ph�   �M$��Q�(x����3҃} �U��}� u!h�j h�   h��j�Lw������u̃}� u3�ݐ���    j h�   h��h\�h��'������   �   �}� tw3�t	�E�   ��E�    �U��U܃}� u!h�j h�   h��j��v������u̃}� u0�]����    j h�   h��h\�h�觉�����   ��-���� "   �"   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���]��������̋�U����} |�}}	�E�   ��E�    �E��E��}� u"h�j jqhp�j�t������u�l���}� u.�%����    j jqhp�h@�h��r���������   �}�t�U���t	�E�    ��E�   �E�E�}� u"h8�j jvhp�j�t������u�'l���}� u+襍���    j jvhp�h@�h8�����������/�}�u�U���N��E���N�M��U�E���N�E���]������������������������������������������������������������������������������������������̋�U����} |�}}	�E�   ��E�    �E�E��}� u%h�j h�   hp�j�s������u�k���}� u0蒌���    j h�   hp�hH�h��܅����������c�}�u�U���N�Q�E���N�M��}�uj��@��U���N�'�}�uj��@��M���N��U�E���N�E���]��������������������������������������������������������������̋�U��Q���E��M���E���]������������������̋�U���]����̋�U��j�h�0h�d�    P���PP  �p����A1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�r����ƅ���� h�  j ������Q�r����3�f������h�  j ������P��q����ƅЯ�� h�  j ��ѯ��Q��q�����} |�}|����*  �E�    �}��   h�N������   j h  hp�h��hP�j
h   ��п��R�EP�,�����P�Y|����h ��ܒ�} t�M�������
ǅ�����������R�ܒh ��ܒ��п��P�ܒhI�ܒ�dh��ǅ���������=  �} ��   ǅ̯��    �ŉ�����ȯ��踉���     �UR�EPh�  h   ��Я��Q�ӆ������̯����̯�� }*j h*  hp�h��h\fj"j�c����R�Vk���� �S�����ȯ�����̯�� }8j h-  hp�h��hH�h<�h   ��Я��R�L�����P�{�����}uV�} tǅ����,��
ǅ�����j h2  hp�h��hH�������Ph   ��п��Q�������P�z����j h4  hp�h��hؼ��Я��Rh   ��п��P�f����P�z�����}u�M���N��t8j h9  hp�h��h��hx�h   ��п��P��e����P�8z����j h:  hp�h��h �hIh   ��п��Q�e����P� z�����} ��   ǅį��    �և����������ɇ���     ��п��P�MQ�URh�h�  h   ������P��p������į����į�� }*j hA  hp�h��h\fj"j�h����Q�[i���� �X������������į�� }8j hD  hp�h��hp�h<�h   ������P�Q�����P� y�����:j hH  hp�h��h����п��Qh   ������R������P��x����ǅ����    ǅ����    j�������Ph   ������Q������R�z}����������j hM  hp�h��h��j"j������P�jh���� ������ t8j hO  hp�h��h�hx�h   ������Q�"�����P�<x�����=,� u�=(� �#  ǅ����    ǅ����    j�m�����E�   �,���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un�(���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j�$z����Ã����� �D  �=� t?ǅ����    ������R������P�MQ������tǅ����   ������������������ ��   �E���N��t>�U�<��N�t1j ������P������Q�/n����P������R�E���NQ����U���N��t������Q�ܒ�U���N��twƅп�� �} t9j h�  hp�h��hP�j
h   ��п��Q�UR�~����P��u������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�d�����������E������   ��}uh�N�(�Ë������M�d�    Y_^[�M�3���c����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h 1h�d�    P���\�  �\f����A1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q��g����3�f������h�  j ������P��g����ƅ���� h�  j ������Q�g����3�f��Џ��h�  j ��ҏ��P�g�����} |�}|����.  �E�    �}��   h�N������   j h�  hp�h��h��j
h   ��Я��Q�UR��u����P�%r����h8����} t�E������
ǅ���������Q��h������Я��R��h�����0^��ǅ���������A  �} ��   ���� ��ȏ������     �MQ�URh�  h   ��Џ��P�x������̏����̏�� }*j h  hp�h��h\fj"j�9���Q�,a���� �)����ȏ�����̏�� }8j h  hp�h��h@�h�h   ��Џ��P������P��p�����}uV�} tǅ�����
ǅ�����j h  hp�h��h������Qh   ��Я��R�{����P�p����j h  hp�h��h����Џ��Ph   ��Я��Q��[����P�[p�����}u�U���N��t8j h  hp�h��hH�h@�h   ��Я��Q�[����P�p����j h  hp�h��h��h��h   ��Я��R�g[����P��o�����} ��   ǅď��    �}��� �������}���     ��Я��Q�UR�EPh��h   h   ������Q��`������ď����ď�� }*j h  hp�h��h\fj"j�>}���R�1_���� �.}�����������ď�� }8j h  hp�h��hx�h�h   ������R��}����P��n�����:j h"  hp�h��h`���Я��Ph   ������Q�}����P�n����ǅ����    j h(  hp�h��h��j"jj�������Rh   ������Pj �N[����P�[^���� ������������ t8j h*  hp�h��h��hx�h   ������Q�X}����P�'n�����=,� u�=(� �#  ǅ����    ǅ����    j�c�����E�   �,���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un�(���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j�p����Ã����� �g  �=� t?ǅ����    ������R������P�MQ������t������������ǅ����   ������ �  �E���N���[  �U�<��N��J  �E���NQ�H�����������t�Jj ������R������P�c����P������Q�U���NP�����t��   �$���t��   ǅ���    j h{  hp�h��hؿj"jj�������Qh   �����R�����P�X����P�[���� ���������� t>�����Pt5j ������Q������R��b������P������P�M���NR����@����� v������������j ������Q�����R�����P�M���NR����E���N��t������R���E���N��ty3�f��Я���} t9j h�  hp�h��h��j
h   ��Я��P�MQ�Qn����P�j������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ�Y�����������E������   ��}uh�N�(�Ë������M�d�    Y_^[�M�3��X����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���@��A3ŉE��E�    �b���E��E�    �E�    �E�    �=�m ��   h�� ��Eԃ}� u3��  h@��E�P����E��}� u3��  �M�Q����mh��U�R���P����mẖ�E�P���P����mh ��M�Q����E��U�R����m�=�m th���E�P���P����m��m;M�th��m;U�t]��mP�ܑ�EЋ�mQ�ܑ�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W��m;M�t��mR�ܑ�Eȃ}� t�UȉE�}� t*��m;E�t ��mQ�ܑ�Eă}� t
�U�R�UĉE䡄mP�ܑ�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��T����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} u3��k  3��} ���E��}� uh0�j j7h��j�AY������u̃}� u0��r���    j j7h��h��h0��l�����   �  �} t�U;U��   �EPj �MQ�Y����3҃} �U��}� uh��j j=h��j�X������u̃}� u-�Hr���    j j=h��h��h���k�����   �~�M;M҃��U�uhP�j j>h��j�VX������u̃}� u-��q��� "   j j>h��h��hP��4k�����"   ��   ��MQ�UR�EP�ab����3���]�������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����������������������̋�U���D�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� u!hoj h�   hh�j��V������u̃}� u1�p���    j h�   hh�hL�ho��i��������Z  3Ƀ} ���M̃}� u!hx�j h�   hh�j�V������u̃}� u1�p���    j h�   hh�hL�hx��hi���������   �E�E��M��AB   �U�E�B�M�U��E��@����M�Qj �UR�E�P�p�����E��} u�E��   �M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj �i�����EċE�H���M��U�E��B�}� |!�M�� 3�%�   �E��M����E���M�Qj ��h�����E��E���]��������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�'f������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ��\������]����������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�`������]������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ��^������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�;\������]��������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�]_������]����������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR��]������]��������������������̋�U��Q�E�E��M�Q�UR�Y������]����������������̋�U��Q�E�E��M�Q�UR�U������]����������������̋�U��Q�E�E��M�Q�UR�EP��T������]������������̋�U��Q�E�E��M�Q�UR�EP�fe������]������������̋�U��Q�} t��}��E�P�V  ���M��} t
��  �U���]��������������������������̋�U�����}��E�P�
  ���E��=�� t�]�M�Q��  ��E���E���]�������������������������������̋�U��QV�}���=�� t�E�P�  �����w  ����M�Q�  ��^��]�������������������������������̋�U����} t^��}��E�P��  ���E�M#M�U��#U�ʉM��E�;E�t'�M�Q�Z  ��f�E��m���}��U�R�  ���E��E�M���} t)�=�� t�UR�EP��  ���M��	�U�    �   ��]��������������������������������������������̋�U��E%����P�MQ��O����]��������������������̋�U�����}��E�P��  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�`  ��f�E��m���}��U�R�  ���E�=�� tB�EP�MQ��  ���E�U�#���E�#��;�t�E�E�   ����E�E����E��]������������������������������������������������̋�U����} 	 u>�}�u8��}��E�%=  ==  u$�=�� t�]��M�����  ���  u�;��7j h[  h��hl�h���U������R�EPj �`����P�Z������]��������������������������������������̋�U�����P��� �E�����E���R	  �}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]�������������������������̋�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]��������������������������������������������������������������������������������������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��������������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�������������������������������������̋�U��Q�!K���E��E�P�)  ����]������������������̋�U��Q�]��e���U��E�P��  ����]��������������̋�U����E%�E�]��M�Q�   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R��  ���E��E�P�/H�����]��M�Q�2   ����]�������������������������������������������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]��������������������������������������������������������������������������������������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]��������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]��������������������������������������������̋�U��Q�E��  �E�P��C������]�������������������̋�U���]����̋�U���]����̋�U����N���E��E��Hp����Ƀ��M��U�U��E����E��}�wC�M��$��d�U��Bp���M��Ap�   �U��Bp����M��Ap�   �   ��H�����u3�t	�E�   ��E�    �E�E�}� u!h�j h�   h��j�:D������u̃}� u.��]���    j h�   h��hh�h��W���������E���]ÐodjdBdVd�����������������������������������������������������������������������̋�U��j�hP1h�d�    P��SVW��A1E�3�P�E�d�    �=LKHJtAj�D�����E�    hHJhLK�Z�����LK�E������   �j��Q����ËM�d�    Y_^[��]�����������������������������������������������̋�U��j�hp1h�d�    P��SVW��A1E�3�P�E�d�    �} ��   j��C�����E�    �E�x t.�M�QR�(���u�E�xhBtj�M�QR��Q�����E������   �j�Q����ËE�8 tcj�{C�����E�   �M�R�W�����E�8 t#�M��: u�E�8HJt�M�R��=�����E������   �j�P����ËE� 𭺋M�A�j�UR�*Q�����M�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��EP�C����]�������������̋�U����E�    �} |�}�} u3��  he  h��jjj��Y�����E��}� u�Z���    3��  hj  h��jjh�   �Y�����M���U��: u j�E�P�P�����<Z���    3��8  hp  h��jjh   �OY�����E��M��U��Q�}� u0j�E��Q��O����j�U�R�O������Y���    3���   hHJ�E��Q�P  ���UR�EP�M��R�z  ����u3�E��Q�gU�����U��P��;����j�M�Q�LO�����E�    �x�U��BP�M���BP�A������tDj�M��QR�O�����E��Q�U�����U��P�m;����j�M�Q��N�����E�    ��U��B�    �M��Q�   �E���]���������������������������������������������������������������������������������������������������������������������������������̋�U��VW�} t0�} t*�E;Et"�u�6   �}�M�    �UR�8S����_^]�������������������������������̋�U��EP�MQ�rJ����]���������̋�U��j�h�1h�d�    P���SVW��A1E�3�P�E�d�    �E�    �3G���E�h�  h��jjj��V�����E�}� u�W���    3��   �N���vP���E�M��Ql��E�M��Qh�Pj��>�����E�    �E�Q�AR�����E������   �j�WL�����j��>�����E�   �U�BP���E������   �j� L����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������̋�U���O��]����̋�U��j�h�1h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �EԉE؃}� u!h��j h&  h��j�]<������u̃}� u0��U���    j h&  h��h��h���8O����3��  �=E���E��LL���U܋Bp���M܉Ap�E�    h1  h��jjh�   ��T�����E�}� �  j�=�����E�   �U܋BlP�M�Q��������E�    �   �j�mJ����Ã}� ��   �UR�EP�M�Q��  ���E��}� ��   �} th�H�UR��>������t
��m   j�<�����E�   �E�P�M܃�lQ��Q�����U�R�P�����E܋Hp��u$��H��u�E܋HlQhLK�Q�����
  �E�    �   �j�I�������U�R�5P�����E�P�6�����E������   ��M܋Qp���E܉PpËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��LK���   � O�LK���   �8O�LK���   ��R]���������������������̋�U���   ��A3ŉE��} tC�} t�EP�MQ�UR�  ����T�����E���M�TH��T�����T����E��|  ǅd���   ǅh���    �} �O  �M���L�'  �E�H��C�  �U�B��_�  �M��`���h���`���R�:0������\�����\��� t"��\���+�`�����X���t��\������;u3���  ǅl���   ���l�������l�����l���N��X���Q��`���R��l���k���x�Q�HJ������u"��l���k���x�P�;����9�X���u�뚋�\�������\���h���\���R�/������X�����X��� u��\������;t3��$  ��l���|j h�  h��h��h@���X���R��\���Ph�   ��p���Q�*5����P�@C������X���Ƅp��� ��p���P��l���Q�UR��  ����t��h�������h�����\����X�����`�����`������t��`�������`�����`�������7�����h��� t�MQ��  ����P����
ǅP���    ��P����U��  �EPj j h�   ��p���Q�UR�L�����E��}� ��   ǅl���    ���l�������l�����l���|��l��� tn��l������U�D
HP��p���Q�:������t;��p���R��l���P�MQ�  ����t��h�������h����
ǅd���    ���h�������h����l�����d��� t�MQ��  ���E��0��h��� t�UR�  ����L����
ǅL���    ��L����E���MQ�  ���E��E��M�3��/����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ��A3ŉE�ǅX���    ǅT���    �=����D�����D����  ��l���ǅH���   �MQ��@���R��L���Ph�   ��p���Q�UR� J������u3��  �E���M�THR��p���P�7������u�M���U�D
H�a  ��p���P�O7��������T���h�  h��j��T���Q��,������X�����X��� u3��  �U���E�LH��8����U�E�L���<���j�Uk��E�L$Q��0���R�=�����E�H��\���j h  h��h��h���p���R��T�����P��X�����Q��M����P��>������X������E���M�TH��L����E�M�T�j��L���R�Ek��M�T$R�)=�����}�
  �E��@����H��H�����l����L���T����(�����,���ǅ`���    ���`�������`�����`���;�H�����   �U��`�����l����R;�uJ��`��� t=��`�����l������D���l�����A��`�����l�����(����Ћ�,����L��]�V��`�����l����ЋT���d�����h�����`�����l�����(�������,����T���d�����(�����h�����,����#�����`���;�H�����   j�E�HQ�U�BP��8���Qjh��jj ��>���� ����   ǅ$���    ���$�������$�����$���s$��$�����E8������  ��$���f��U8�����h�   ��NP��8���Q�_;������u��l����B   ���l����@    ���l����A    ��l����E�H�
�U��l����H���   �}u�U��@����B�MQ�Uk������Ѓ���tG�M���U��8����D
Hj��X���Q��?�����U�E��<����L��U��\����B3��   ��8����Ht{�M���U�D
PP�(���uc3�uj j h[  h��j�0������u�j�E���M�TPR�Y?����j�E���M�TTR�A?�����E���M�DL    ��X��� t��X����   �E���M��X����TP�E���M�DH�M�3��)����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�    �E�    �E�    �E�U  ht  h��j�E�P�$'�����E�}� u3��  �M���M��U���U��E��  �M��   �E�   �	�U����U��E����M�THRh���E�k���x�Qj�U�R�E�P�B%�����}�}kj h�  h��h �h��h��M�Q�U�R�v$����P��8�����E������M�THR�E����M�THR�0������t�E�    �  �}� ��   �E�xP tD�M�QPR�(���u33�uj j h�  h��j��,������u�j�U�BPP�<�����M�yT tD�U�BTP�(���u33�uj j h�  h��j�s,������u�j�E�HTQ��;�����U�BT    �E�@L    �M�U�QP�E�M��HH�E���   ��   j�U�R�;�����E�xP tD�M�QPR�(���u33�uj j h�  h��j��+������u�j�U�BPP�A;�����M�yT tD�U�BTP�(���u33�uj j h�  h��j�+������u�j�E�HTQ��:�����U�BT    �E�@L    �M�AP    �U�BH    �E�@h�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����   ��A3ŉE��3���   �E�E��(�E��M�� �M�U��,�U��E�   �E��   �E��E��   �E�    �} u3��-  �} t�} u3��  �M���Cuv�E�H��ukj h�  h��h��h0�h,��UR�EP�D����P�l5�����} t3ɋUf�
3��Mf�A3ҋEf�P�} t	�M�    �E�  �UR��,�����E��}��   s0�EP�M�Q�-�������  �UR�E�P��,��������   ǅ@���    ǅD���    �MQ��H���R�*������t3��  ��H���P�M�Q��H���R��+������u3���   �E��H�U��
��H���P�M�Q�U�R�p-�����E���t�}��   s�U��@����E���D����
ǅ@����Kj h�  h��h��h����D�����Q��@���R�E�P�M�Q��%����P�4�����} tj�U�R�EP�2�����} tj�M�Q�UR�~2����j h  h��h��h0��E�P�MQ�UR��B����P�3�����E��M�3���!����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�]�������̋�U����E�E��E�    �	�M����M��U�;U}A�E����E�j h  h��h\�h���M��Q�R�EP�MQ������P�l2������E�    ��]��������������������������������������������̋�U���h�   j �EP�'�����M���u3���  �E���.uX�U�B��tMj h*  h��hX�hX�j�M��Qj�U�   R�#����P�1�����Eƀ�    3��e  �E�    �	�M����M�hT��UR�������E��}� u����1  �EE���M��}� uI�}�@sC�U���.t:j h8  h��hX�h`��E�P�MQj@�UR�#����P�1�����   �}�uI�}�@sC�E���_t:j h;  h��hX�hp��M�Q�URj@�E��@P�"����P��0�����_�}�uT�}�sN�M���t	�U���,u=j h>  h��hX�hx��E�P�MQj�U�   R�Y"����P�o0���������)�E���,u��M���u��U��E�L�M����3���]����������������������������������������������������������������������������������������������������������������������������������������̋�U��j hT  h��h�h���EP�MQ�UR�>����P�{/�����E�H@��t�U��@Rh|�j�EP�MQ�p�����U���   ��t!�M���   Qhx�j�UR�EP�A����]����������������������������������������������̋�U����EP�M��.���M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M��f"��P�.   ��$�E�M��F=���E��]�������������������������̋�U��� �} ~,�EP�MQ�%  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R���E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R�%����P�78�����E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R����u
�Y  �T  j j �E�P�M�Q�UR�EP���E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR����u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�~$����P�07�����E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ����u�V�T�}  u+j j j j �U�R�E�Pj �M$Q���E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P���E��}� t�M�Q�8�����U�R�8�����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U����EP�M���)���M��v����U���   �P�� �  �M�M��I9���E��]����������������������������̋�U��j �EP�4 ����]�����������̋�U��h  �EP�*����]�������̋�U��h  �EP��)����]�������̋�U��j�EP��)����]����������̋�U��j�EP�)����]����������̋�U��j�EP�)����]����������̋�U��j�EP�x)����]����������̋�U��j�EP�X)����]����������̋�U��j�EP�8)����]����������̋�U��h�   �EP�)����]�������̋�U��h�   �EP��(����]�������̋�U��j�EP��(����]����������̋�U��j�EP�(����]����������̋�U��j�EP�(����]����������̋�U��j�EP�x(����]����������̋�U��h  �EP�U(����]�������̋�U��h  �EP�5(����]�������̋�U��hW  �EP�(����]�������̋�U��hW  �EP��'����]�������̋�U��h  �EP��'����]�������̋�U��h  �EP�'����]�������̋�U��j �EP�'����]����������̋�U��j �EP�x'����]����������̋�U���E=�   ���]������������̋�U��Qh  �EP�4'������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP��&������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�&������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�D&������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ����������������������������XY�$�����������XY�$�����������XY�$����������̋�U���SVWd�5    �u��E��j �EP�M�Q�UR��%���E�H����U�Jd�=    �]��;d�    _^[��]� ����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�g-���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�-���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ��,���� �E�_^[�E���]��������������������̋�U��E�HQ�U�B(Pj �M�QR�����]� �����������������������̋�U����E�    �E����A�M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ�n���E�E�d�    �E��]����������������������������������̋�U��Q��E�H3M����j �MQ�U�BP�M�QRj �EP�M�QR�EP�+���� �E��E���]��������������������̋�U���8S�}#  u�.��M��   ��   �E�    �Eܠ���A�M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M�� �����   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]��������������������������������������������������������������������̋�U��QS��E�H3M�=���M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ��)���� �U�z$ u�EP�MQ� *��j j j j j �U�Rh#  ������E��]�c�k ��   [��]���������������������������������������������������̋�U��Q�} �E�HSV�pW�M�����|8����u�����E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v����M�_��^��[��]��������������������������������̋�U��EV�u��������   �N�������   ��^]��������������������̋�U��������   ��t�M9t�@��u��   ]�3�]�������������������̋�U��V�f���u;��   u�V���N���   ^]��E�����   �x t�H;�t���x u�^]����V�P^]�������������������������̋�U����EP�M�����M$Q�U R�EP�MQ�UR�EP�MQ�M��
��P�2   �� �E�M���-���E��]�����������������������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP���E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP�k����P�)�����E���E�    �M�M��}� u3��a�U���Rj �E�P�g�����M�Q�U�R�EP�MQj�UR���E��}� t�EP�M�Q�U�R�EP���E��M�Q�*�����E���]�����������������������������������������������������������������������̋�U��Q�E�x  toj?h��jhd  j��*�����E��}� u
�   �   �MQ�U�R��   ����t!�E�P�X*����j�M�Q�+!�����   �}�U�ǂ�      ��E��H�E���   �HtJ�M���   �´   R�(���u0�E���   ���    h��j jOh(�j�H������u̋E�M����   3���]����������������������������������������������������������������̋�U����E�    �E�HB�M��U�BD�E��} u�����  �M�M��E�    �U��Rj1�E�Pj�M�Q������E�E�U��Rj2�E�Pj�M�Q������E�E�U��Rj3�E�Pj�M�Q�����E�E�U��Rj4�E�Pj�M�Q�����E�E�U��Rj5�E�Pj�M�Q�d����E�E�U��Rj6�E�Pj�M�Q�C����E�E�URj7�E�Pj�M�Q�%����E�E�U�� Rj*�E�Pj�M�Q�����E�E�U��$Rj+�E�Pj�M�Q������E�E�U��(Rj,�E�Pj�M�Q������E�E�U��,Rj-�E�Pj�M�Q�����E�E�U��0Rj.�E�Pj�M�Q�����E�E�U��4Rj/�E�Pj�M�Q�_����E�E�U��Rj0�E�Pj�M�Q�>����E�E�U��8RjD�E�Pj�M�Q�����E�E�U��<RjE�E�Pj�M�Q������E�E�U��@RjF�E�Pj�M�Q������E�E�U��DRjG�E�Pj�M�Q�����E�E�U��HRjH�E�Pj�M�Q�����E�E�U��LRjI�E�Pj�M�Q�x����E�E�U��PRjJ�E�Pj�M�Q�W����E�E�U��TRjK�E�Pj�M�Q�6����E�E�U��XRjL�E�Pj�M�Q�����E�E�U��\RjM�E�Pj�M�Q������E�E�U��`RjN�E�Pj�M�Q������E�E�U��dRjO�E�Pj�M�Q�����E�E�U��hRj8�E�Pj�M�Q�����E�E�U��lRj9�E�Pj�M�Q�p����E�E�U��pRj:�E�Pj�M�Q�O����E�E�U��tRj;�E�Pj�M�Q�.����E�E�U��xRj<�E�Pj�M�Q�����E�E�U��|Rj=�E�Pj�M�Q������E�E�U�   Rj>�E�Pj�M�Q������E�E�U�   Rj?�E�Pj�M�Q�����E�E�U�   Rj@�E�Pj�M�Q�����E�E�U�   RjA�E�Pj�M�Q�\����E�E�U�   RjB�E�Pj�M�Q�8����E�E�U�   RjC�E�Pj�M�Q�����E�E�U�   Rj(�E�Pj�M�Q������E�E�U�   Rj)�E�Pj�M�Q������E�E�U�    Rj�E�Pj�M�Q�����E�E�U�¤   Rj �E�Pj�M�Q�����E�E�U�¨   Rh  �E�Pj�M�Q�]����E�E�U�°   Rh	  �E�Pj �M�Q�6����E�E�U�E����   �M���   Qj1�U�Rj�E�P�����E�E�M���   Qj2�U�Rj�E�P������E�E�M���   Qj3�U�Rj�E�P�����E�E�M���   Qj4�U�Rj�E�P�����E�E�M���   Qj5�U�Rj�E�P�v����E�E�M���   Qj6�U�Rj�E�P�R����E�E�M���   Qj7�U�Rj�E�P�.����E�E�M���   Qj*�U�Rj�E�P�
����E�E�M���   Qj+�U�Rj�E�P������E�E�M���   Qj,�U�Rj�E�P������E�E�M���   Qj-�U�Rj�E�P�����E�E�M���   Qj.�U�Rj�E�P�z����E�E�M���   Qj/�U�Rj�E�P�V����E�E�M���   Qj0�U�Rj�E�P�2����E�E�M���   QjD�U�Rj�E�P�����E�E�M���   QjE�U�Rj�E�P������E�E�M���   QjF�U�Rj�E�P������E�E�M���   QjG�U�Rj�E�P�����E�E�M��   QjH�U�Rj�E�P�~����E�E�M��  QjI�U�Rj�E�P�Z����E�E�M��  QjJ�U�Rj�E�P�6����E�E�M��  QjK�U�Rj�E�P�����E�E�M��  QjL�U�Rj�E�P������E�E�M��  QjM�U�Rj�E�P������E�E�M��  QjN�U�Rj�E�P�����E�E�M��  QjO�U�Rj�E�P�����E�E�M��   Qj8�U�Rj�E�P�^����E�E�M��$  Qj9�U�Rj�E�P�:����E�E�M��(  Qj:�U�Rj�E�P�����E�E�M��,  Qj;�U�Rj�E�P��
����E�E�M��0  Qj<�U�Rj�E�P��
����E�E�M��4  Qj=�U�Rj�E�P�
����E�E�M��8  Qj>�U�Rj�E�P�
����E�E�M��<  Qj?�U�Rj�E�P�b
����E�E�M��@  Qj@�U�Rj�E�P�>
����E�E�M��D  QjA�U�Rj�E�P�
����E�E�M��H  QjB�U�Rj�E�P��	����E�E�M��L  QjC�U�Rj�E�P��	����E�E�M��P  Qj(�U�Rj�E�P�	����E�E�M��T  Qj)�U�Rj�E�P�	����E�E�M��X  Qj�U�Rj�E�P�f	����E�E�M��\  Qj �U�Rj�E�P�B	����E�E�M��`  Qh  �U�Rj�E�P�	����E�E�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u�W  j�E�HQ�����j�U�BP������j�M�QR������j�E�HQ������j�U�BP�����j�M�QR�����j�E�Q�����j�U�B P�����j�M�Q$R�{����j�E�H(Q�j����j�U�B,P�Y����j�M�Q0R�H����j�E�H4Q�7����j�U�BP�&����j�M�Q8R�����j�E�H<Q�����j�U�B@P������j�M�QDR������j�E�HHQ������j�U�BLP������j�M�QPR�����j�E�HTQ�����j�U�BXP�����j�M�Q\R�|����j�E�H`Q�k����j�U�BdP�Z����j�M�QhR�I����j�E�HlQ�8����j�U�BpP�'����j�M�QtR�����j�E�HxQ�����j�U�B|P������j�M���   R������j�E���   Q������j�U���   P�����j�M���   R�����j�E���   Q�����j�U���   P�|����j�M���   R�h����j�E���   Q�T����j�U���   P�@����j�M���   R�,����j�E���   Q�����j�U���   P�����j�M���   R������j�E���   Q������j�U���   P������j�M���   R�����j�E���   Q�����j�U���   P�����j�M���   R�x����j�E���   Q�d����j�U���   P�P����j�M���   R�<����j�E���   Q�(����j�U���   P�����j�M���   R� ����j�E���   Q������j�U���   P������j�M���   R������j�E���   Q�����j�U��   P�����j�M��  R�����j�E��  Q�t����j�U��  P�`����j�M��  R�L����j�E��  Q�8����j�U��  P�$����j�M��  R�����j�E��   Q������j�U��$  P������j�M��(  R������j�E��,  Q������j�U��0  P�����j�M��4  R�����j�E��8  Q�����j�U��<  P�p����j�M��@  R�\����j�E��D  Q�H����j�U��H  P�4����j�M��L  R� ����j�E��P  Q�����j�U��T  P��
����j�M��X  R��
����j�E��\  Q��
����j�U��`  P�
����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �E�    �E�E��E�    �M�y u�U�z �  jeh��jjPj�-�����E�}� u
�   ��  �E���   �   �}��jqh��jj�U������E�}� uj�M�Q�s�����   �z  �U��    �E�x �:  j}h��jj�������E��}� u&j�M�Q�)����j�U�R������   �"  �E��     �M�Q>�U��E�Pj�M�Qj�U�R�������E�E�E��Pj�M�Qj�U�R������E�E�E��Pj�M�Qj�U�R������E�E�E��0Pj�M�Qj�U�R�a�����E�E�E��4Pj�M�Qj�U�R�@�����E�E�t0�E�P�����j�M�Q�@����j�U�R�2��������;  �E�HQ�  ���@�E�    �U��N��M��N�Q�E��N�H�U� O�B0�M�O�Q4�E��    �}� t	�M��   ��E�    �E�    �E��N�U���    tA�E���   Q�(���u-�U���    w!h��j h�   h0�j���������u̋M���    t<�U���   P�(���u(j�M���   R�)����j�E���   Q������U�E����   �M�U쉑�   �E�M䉈�   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�   �E�;�Ntj�U�P�F�����M�Q;�Ntj�E�HQ�'�����U�B;�Ntj�M�QR������E�H0; Otj�U�B0P�������M�Q4;Otj�E�H4Q������]�����������������������������������������������������̋�U���VW�E�    �E�E��E�    �M�y u�U�z �W  jSh��jjPj������E�}� u
�   ��  jYh��jj��������E��}� uj�E�P������   ��  �M��    �U�z �d  jeh��jj�������E�}� u&j�E�P������j�M�Q������   �s  �U��    �E�H8�M��E�    �U��Rj�E�Pj�M�Q�T�����E�E�U��Rj�E�Pj�M�Q�3�����E�E�U��Rj�E�Pj�M�Q������E�E�U��Rj�E�Pj�M�Q�������E�E�U��Rj�E�Pj�M�Q�������E�E�U�� RjP�E�Pj�M�Q������E�E�U��$RjQ�E�Pj�M�Q������E�E�U��(Rj�E�Pj �M�Q�m�����E�E�U��)Rj�E�Pj �M�Q�L�����E�E�U��*RjT�E�Pj �M�Q�+�����E�E�U��+RjU�E�Pj �M�Q�
�����E�E�U��,RjV�E�Pj �M�Q�������E�E�U��-RjW�E�Pj �M�Q�������E�E�U��.RjR�E�Pj �M�Q������E�E�U��/RjS�E�Pj �M�Q������E�E�U��8Rj�E�Pj�M�Q�e�����E�E�U��<Rj�E�Pj�M�Q�D�����E�E�U��@Rj�E�Pj�M�Q�#�����E�E�U��DRj�E�Pj�M�Q������E�E�U��HRjP�E�Pj�M�Q�������E�E�U��LRjQ�E�Pj�M�Q�������E�E�t@�U�R�e����j�E�P�������j�M�Q������j�U�R�������   �b  �E�HQ�  ����   ��N�}��U���   �M���E���   �U�A�B�M���   �E�J�H�U���   �M�P0�Q0�E���   �U�A4�B4�M��   �}� t	�U��   ��E�    �E�    �E��N�E���    tA�M���   R�(���u-�E���    w!h��j h�   h0�j�9�������u̋U���    t<�E���   Q�(���u(j�U���   P�r�����j�M���   R�^������E�M䉈�   �U�E����   �M�U艑�   3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�  �E�H;�Ntj�U�BP�������M�Q;�Ntj�E�HQ��������U�B;�Ntj�M�QR��������E�H;�Ntj�U�BP�������M�Q;�Ntj�E�HQ�������U�B ;�Ntj�M�Q R�i������E�H$;�Ntj�U�B$P�J������M�Q8;Otj�E�H8Q�+������U�B<;Otj�M�Q<R�������E�H@;Otj�U�B@P��������M�QD;Otj�E�HDQ��������U�BH;Otj�M�QHR�������E�HL;Otj�U�BLP������]�����������������������������������������������������������������������������������������������������������̋�U���������E��E��Hl�M��U�;LKt�E��Hp#�Hu�����E�� O��]�����������������������������̋�U��<O]����̋�U����T����E��E��Hl�M��U�;LKt�E��Hp#�Hu�A����E��U����   ��]�������������������������̋�U��hDO�EP�MQ�t����]��������������������̋�U���<��A3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q�������t	�E�    ��U�R�������E�   �Z  �E�P�M�Q�'������U�U؋E�HQ�U�R�n�������t	�E���E�M�U�A+B9E�}�M�Q�#������E�    �E�   ��   �U�E�;Bk�M�Q�U�R�������E؉E�M�Q+U�UċE�P�M�Q��������U�BP�M�Q��������U�B��P�M�Q�������E�    �E�   �~�U�E�;|B�M�Q�������U܁�   ��U܋E�HQ�U�R�R������E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�������E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3��Y�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ��������u�U�R�EP�m������E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������������������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]��������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P�������E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R��������E��ȋE���]������������������������������������������������������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]����������������̋�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]����������������������������������̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�����������������������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]������������������������������������������������������������������̋�U��h\O�EP�MQ�$�����]��������������������̋�U�����A3ŉE��E�    �E�H
���  f�M��U�B
% �  f�E�M�Q�U�E�H�M�U����E�j@�M�Q�w�������t�E�   �f�U�f��f�U��E�=�  u�E�   �M�U�Q�E�M��U��E�ЋMf�Q�E��M�3�������]��������������������������������������������������������������̋�U���   ��A3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h��j h�   h��j���������u̃}� u0�V����    j h�   h��h��h��������3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$�4��U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p�����t��$�d��E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h��������$����E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�������$����E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�2������}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�>�����f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3��������]Ë�����U�����������f��$���.��%�@�  ���}���  �{�r���  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����A3ŉE�� S��`�E��} u�   �} }�M�ىM��T��`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP������눋M�3��2�����]�����������������������������������������������������������̋�U���L��A3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�K������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q�!�����f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R������f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]������������������������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]���������������������������̋�U�����A3ŉE��EPj j j �MQ�UR�EP�M�Q�m����� �E�UR�E�P�^������E��}�u	�M���M�E�M�3�������]��������������������������������������̋�U���x��A3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|hX�h<�h��h��j�U��R�������P�������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   hX�h<�h��h|�j�U��R�w�����P�F������E�@�E�    �   �}�   �uK�}� uEj h�   hX�h<�h(�h�j�M��Q� �����P��������U�B�E�    �Cj h�   hX�h<�h��h��j�E��P�������P�������M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q��������U����?  |f�E�f��f�E��M�Q�U�R�z������Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�`�������}� },�E���%�   �E��	�M����M��}� ~�U�R�n�������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P��������M�Q��������U�R�E�P�
������M�Q��������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3��¿����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�R�E�Q�������E��}� t0�U��Rj�E�HQ�������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�f������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR�1�������]��������������������������������������������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y��������������������������������������������������������������������������������̋�U��j
j �EP������]���������̋�U��EPj
j �MQ�<�����]���������������������̋�U��EP�������]�������������̋�U��EP�MQ�0�����]���������̋�U��j
j �EP�|�����]���������̋�U��EPj
j �MQ�D�����]����������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� �������������������������������������������U��SVWUj j h���u����]_^[��]ËL$�A   �   t2�D$�H�3��ӹ��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h �d�5    ��A3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y �u�Q�R9Qu�   �SQ��O�SQ��O�L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������������������̋�U���8�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uhoj jph�nj�*�������u̃}� u.�����    j jph�nh��ho����������   3Ƀ} ���MЃ}� uhx�j juh�nj�ƽ������u̃}� u.�W����    j juh�nh��hx�����������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P�������E��} u�E��Q�M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �`������EȋE���]������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR������]�������������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!hoj h�  h�nj���������u̃}� u.�����    j h�  h�nh�ho�����������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh��������]������������������̋�U��EP�MQ�URh���{�����]����������������̋�U��EPj �MQhù�M�����]������������������̋�U��EP�MQ�URhù������]����������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uhoj jph�nj�*�������u̃}� u.�����    j jph�nh0�ho����������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh0nj jsh�nj谹������u̃}� u.�A����    j jsh�nh0�h0n�����������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �3������Eă}��t�E���UU�B� �E��x }�����������]��������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh���W������E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh����������E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�j h�   h�nj�$�������u̃}� u1�����    j h�   h�nh��h�������������  �} t�} v	�E�   ��E�    �U�U�}� u!h��j h�   h�nj褶������u̃}� u1�5����    j h�   h�nh��h������������d  �MQ�UR�EP�MQ�URh�褲�����E��}� }U�E�  �}�tI�}���t@�}v:�M��9�As��A�U��	�E���E�M�Qh�   �U��R藶�����}��uu3�t	�E�   ��E�    �M�M��}� u!h\�j h�   h�nj觵������u̃}� u.�8���� "   j h�   h�nh��h\�����������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9�As
��A�E���M����U+щU��E�Ph�   �M��U�D
P赵�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP������]���������������̋�U���,�E������E�    3��} ���E�}� u!h�j h  h�nj��������u̃}� u1�~����    j h  h�nh4�h������������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!h��j h  h�nj�T�������u̃}� u1������    j h  h�nh4�h���/���������|  �M;M��   ������U��EP�MQ�UR�E��P�MQh��;������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9�As��A�U���E���M+ȉM�U�Rh�   �E�M�TR�!����������8"u
�����M������  �`�������U��EP�MQ�UR�EP�MQh�臮�����E��UU�B� �}��u"�}�u�����8"u
�����M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U��E�Ph�   �M��Q�D������}��uu3�t	�E�   ��E�    �E܉E�}� u!h\�j hB  h�nj�T�������u̃}� u.������ "   j hB  h�nh4�h\��/�������������z�}�t\�}���tS�U���;UsH�E����M+�9�As��A�U���E����M+ȉM؋U�Rh�   �E��M�TR�b������}� }	�E�������E��EԋEԋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ������]�����������̋�U����EPj �MQ�UR�EPhù跫�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhù�U������E��}� }	�E�������U��U��E���]������������������������̋�U��j�h2h�d�    P���SVW��A1E�3�P�E�d�    �E������E������}�u!艵���     ����� 	   ��������  �} |�E;<�s	�E�   ��E�    �MԉM܃}� uh��j jMhX�j��������u̃}� u<�����     ����� 	   j jMhX�h@�h����������������C  �E���M���������D
������؉E�uh�j jNhX�j苭������u̃}� u<莴���     ����� 	   j jNhX�h@�h��^������������   �UR萩�����E�    �E���M���������D
��t �MQ�UR�EP�MQ�������E��U��F����� 	   ������     �E������E�����3�uhX�j jYhX�j谬������u��E������   ��MQ������ËE��U�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��UR迶�����E�}��u;�T���� 	   3�u!hX�j h�   hX�j荫������u̃������   �UR�E�P�M�Q�U�R���E��}��u#�$��E��}� t�E�P�D������������>�M���U���������L����U���E���������L�E��U���]������������������������������������������������������������������������̋�U��j�h02h�d�    P���SVW��A1E�3�P�E�d�    �}�u臱���     �
���� 	   ����  �} |�E;<�s	�E�   ��E�    �M؉M��}� uh��j jChP�j��������u̃}� u9�����     ����� 	   j jChP�h@�h������������/  �E���M���������D
������؉E�uh�j jDhP�j菩������u̃}� u9蒰���     ����� 	   j jDhP�h@�h��b���������   �UR藥�����E�    �E���M���������D
��t�MQ�UR�EP�*������E��?����� 	   �����     �E�����3�uhX�j jOhP�j�Ũ������u��E������   ��EP������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U�츐<  �¦����A3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uhP�j jmhP�j蕧������u̃}� u9蘮���     �����    j jmhP�h,�hP��h���������
  �E���M���������D
$�����E��M���t	�U���uo�E��������E�uh�j juhP�j��������u̃}� u9������     �y����    j juhP�h,�h��ƹ���������	  �U���E���������T�� tjj j �EP�l������MQ�C�������td�U���E���������T��   tA�e����EԋEԋHl3҃y �U�E�P�M���U���������Q����E�}� ��  �}� t�U�����  ����E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M���������|
8 ��   �E���M���������D
4P�-�������u!h��j h�   hP�j�?�������u̋U���E���������T4�U��EЊ�M��U���E���������D8    j�U�R�E�P�5��������u�  �   �M��R蕞��������   �E�+E�M+ȃ�v'j�U�R�E�P���������u�O  �MЃ��M��K�U���E���������UЊ�T4�E���M���������D
8   �E����E���  �j�M�Q�U�R�y��������u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R���Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M���������
P�����t�M�+MM�M��U�;U�}�  ��$��E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M���������
P�����t!�M�;M�}�   �U���U�E����E���$��E��   �   �M���t	�U���u{�E�P���������U�;�u�E����E���$��E��R�}� tG�E�   �   f�M��U�R�ѻ�������M�;�u�U����U��E���E���$��E���t�����  �M���U���������L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E���������R�����t �E�E��E�������������+�9M�}���$��E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U���������Q�����t �U�U��U�������������+�9E�}���$��E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  ����t�����t��� u�$��E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E���������R�����t��p���E���p�����$��E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U���������Q�����t�E�    �U��U��	�$��E�}� ��   �}� t0�}�u����� 	   �P����M���U�R�+���������V�L�E���M���������D
��@t�M���u3��%�莶���    ������     ������E�+E�M�3��ǖ����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} uh`�j j.h��j�ʙ������u̋�m����m�U�U�j:ht�jh   �ג�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������������������������������������������������������̋�U����}�u����� 	   3��   �} |�E;<�s	�E�   ��E�    �M��M��}� uh��j j(h@�j苘������u̃}� u*����� 	   j j(h@�h(�h���i�����3���E���M���������D
��@��]���������������������������������������������������̋�U�츘O]����̋�U��Q�= � u� �   ��= �}
� �   h�   h��jj� �P胰������m�=�m u?� �   h�   h��jj� �Q�N�������m�=�m u
�   �   �E�    �	�U����U��}�}�E����O�M���m�����E�    �	�E����E��}�}f�M����U����������<�t8�M����U����������<�t�M����U����������< u�M���ǁ�O�����3���]������������������������������������������������������������������������������������̋�U���6�����]��t�o���j��mQ蘥����]�������������������̋�U��}�Or4�}�Qw+�E-�O����P�,������M�Q�� �  �E�P��M�� Q���]�������������������������������̋�U��}}#�E��P�Ж�����M�Q�� �  �E�P��M�� Q���]�������������������̋�U��}�Or4�}�Qw+�E�H������U�J�E-�O����P��������M�� Q���]�������������������������������̋�U��}}#�E�H������U�J�E��P臣������M�� Q���]�������������������̋�U��Q3��} ���E��}� uh��j j)h �j�`�������u̃}� u+�����    j j)h �h��h���>����������U�B��]�������������������������������̋�U��j�hP2h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E؃}� uhoj j6h��j褓������u̃}� u.�5����    j j6h��ht�ho肦��������   �U�U������� Pj蕋�����E�    �Р���� P輒�����E܋E�Pj �MQ負���� P�۠�����E�螠���� P�U�R�������E������   ��{����� Pj�g�����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP��������]������������̋�U��Q�E�E��M�Q�UR�EP��������]������������̋�U��Q�E�E��M�Qj �UR��������]��������������̋�U��Q�E�E��M�Q�UR�EP�ɗ������]������������̋�U��Q�E�E��M�Qj �UR蛗������]��������������̋�U�����A��3�9�m���M��} t��A���U���E�    �E���m�E���]������������������������̋�U�졐A��3�9�m����]��������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh��j jJh�j荐������u̃}� u0�����    j jJh�h��h���k������   �\  �UR�M��(����M�蟏��� �x ��   �M���   ~C�} t�} v�URj �EP趐����褩��� *   虩����M؍M��@����E���  �} tw3�;U��؉E�uh�Mj j]h�j趏������u̃}� u=�G���� "   j j]h�h��h�M蔢�����E�"   �M��˩���E��x  �U�E��} t	�M�   �E�    �M�蝩���E��J  �=  �E�    �U�Rj �EP�MQj�URj �M��w���� �HQ���E��}� t
�}� ��   �}� ��   �$���z��   �} t�} v�URj �EP�n�����3�t	�E�   ��E�    �U��U܃}� uh\�j j{h�j臎������u̃}� u:����� "   j j{h�h��h\��e������E�"   �M�蜨���E��L�ާ��� *   �ӧ����MȍM��z����E��*�} t�U�E���E�    �M��X����E���M��K�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�?�����]��������������̋�U��� �E������EP�M��ȗ���M��?���P�MQ�M��1�������   P�MQ�U�R�������E�}� u�E��E���E������M��M�M������E��]�����������������������������������������̋�U����E�����j �EP�D���P�MQ�U�R�c������E��}� u�E��E���E������E��]���������������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uhp�j jEh��j蠋������u̃}� u.�1����    j jEh��h��hp��~���������  �MQ�M��=����} �  �M�誊����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M��c����E��O  �M����M��U���U뱋E��EԍM��9����E��%  �  �MQ�URj��EPj	�M�� �����QR���E��}� t�E����EЍM������E���  �$���zt*�"���� *   3ɋUf�
�E������M�蹤���E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M�脉��P�M��R艋������t@�E��H��u,蠣��� *   3ҋEf��E������M��7����E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M�������QR���E��}� u*�.���� *   3��Mf��E������M��ţ���E��   �U��U��M�诣���E��   �   �M�覈��� �x u�MQ襌�����E��M��{����E��j�`j j j��URj	�M��l���� �HQ���E��}� u!蒢��� *   �E������M��1����E�� ��U����U��M������E���M�������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�UR�EP�u�����]�����������������̋�U��=�m uhPK�EP�MQ�UR��������j �EP�MQ�UR������]�����������������������������̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!h�j h�   h��j��������u̃}� u3�s����    j h�   h��h��h�轙�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���E��M���Qh�   �U��R�������} t	�E�     �MQ�M������U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h��j h  h��j���������u̃}� u@�q����    j h  h��h��h��軘�����E�   �M������E���  �M�����P�E�P�MQ�UR�9������E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���M��U���Rh�   �E��P迅����譞����MЍM��T����E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9�As��A�M��	�U���U��E���Ph�   �M��Q�#������U�9U����E�u!h��j h  h��j�I�������u̃}� u=�ڝ��� "   j h  h��h��h���$������E�"   �M��[����E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM�� ����Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�j jh�j�h�������u̃}� u0������    j jh�h��h��F������   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U��E�Ph�   �M��Q�|�����3҃} �U��}� uhD�j jh�j裁������u̃}� u0�4����    j jh�h��hD�联�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9�As
��A�E��	�M���M܋U�Rh�   �E��P舁���������t3�t	�E�   ��E�    �E؉E�}� uh(�j j h�j蘀������u̃}� u0�)����    j j h�h��h(��v������   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9�As
��A�E��	�M���MԋU�Rh�   �E��P�z���������t3�t	�E�   ��E�    �EЉE�}� uh̘j j*h�j�������u̃}� u-����� "   j j*h�h��h̘�h������"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9�As��A�U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR�����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uh�Nj jfh��j�>}������u̃}� u0�ϖ���    j jfh��h��h�N�������   ��  3�;U��؉E�uh��j jgh��j��|������u̃}� u0�m����    j jgh��h��h��躏�����   �  �U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���UԋE�Ph�   �M��Q��|����3҃} ��;U��؉E�uhP�j jih��j�|������u̃}� u0謕��� "   j jih��h��hP���������"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uh�j jjh��j�{������u̃}� u0�0����    j jjh��h��h��}������   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!h��j h�   h��j�z������u̃}� u0�&���� "   j h�   h��h��h���p������"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ������]�����������������̋�U��j �EP�MQ�UR�EP�T���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!h�Nj h>  h��j�x������u̃}� u3覑���    j h>  h��hX�h�N��������   �,  3�;U���؉E�u!h��j h?  h��j�w������u̃}� u3�>����    j h?  h��hX�h��舊�����   ��  �U�� �}��tI�}����t@�}�v:�EЃ�9�As��A�M��	�UЃ��ŰE�Ph�   �Mԃ�Q��w����3҃} ��;U���؉E�u!hP�j hA  h��j��v������u̃}� u3�w���� "   j hA  h��hX�hP���������"   ��  �}r�}$w	�E�   ��E�    �UȉU܃}� u!h�j hB  h��j�dv������u̃}� u3������    j hB  h��hX�h��?������   �{  �E�    �MԉM��} t+�U��-�E����E��M����M��U�ڋE�� �؉U�E�M��M�U3�PR�MQ�UR谏���E�E3�QP�UR�EP�����E�U�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} w�} v�U�;U�r��E�;E�rl�M�� �U�;U���؉E�u!h��j hf  h��j�+u������u̃}� u0輎��� "   j hf  h��hX�h���������"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�B���]����������������̋�U���x��A3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uh�j jfh��j�#s������u̃}� u.贌���    j jfh��hp�h�����������8  �UR�M���}���} �.  �M��-r��� �x ��   �M�;Msp�U�=�   ~"�G���� *   �E������M������E���  �MM��U���M��E���E��u�M��M��M�谌���E��  �U����U�눋E��E��M�菌���E��  �  �M��q������   ��   �} v�UR�EP�  ���E�M�Qj �UR�EP�MQ�URj �M��>q��� �HQ���E��}� t3�}� u-�UU��B���u	�M����M��U��U��M������E���  �1���� *   �E������M��Ћ���E���  ��  �E�Pj �MQ�URj��EPj �M��p����QR���E��}� t�}� u�E����E��M��y����E��j  �}� u�$���zt"觊��� *   �E������M��F����E��7  �M�;M�  �U�Rj �M��0p��� ���   Q�U�Rj�EPj �M��p����QR���E�}� t�}� t"�3���� *   �E������M��Ҋ���E���  �}� |�}�v"����� *   �E������M�褊���E��  �E�E�;Ev�M��M��M�胊���E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M��.����E��  벋U���U������E��E��M������E���   ��   �M���n����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"����� *   �E������M�衉���E��   �Ũ��U�벋ẺE��M�耉���E��t�j�M�Qj j j j��URj �M��kn��� �HQ���E��}� t�}� t苈��� *   �E������M��*����E���U����U��M������E���M������M�3��h����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�������������������������������������̋�U��EP�MQ�UR�EP������]�����������������̋�U��j �EP�MQ�UR������]�������������������̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h��j h@  h��j�"l������u̃}� u3賅���    j h@  h��hl�h����~�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U��E�Ph�   �M��Q�7l�����} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h��j hL  h��j�0k������u̃}� u3������    j hL  h��hl�h���~�����   �  �MQ�U�R�EP�MQ�(������E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9�As��A�M��	�U���U؋E�Ph�   �M��Q�$k��������� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9�As
��A�E��	�M���MԋU�Rh�   �E��P�j�����M9M���ډU�u!h8�j hd  h��j��i������u̃}� u0�S���� "   j hd  h��hl�h8��|�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�h����]�����������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!hoj h�   hh�j�h������u̃}� u1蘁���    j h�   hh�h8�ho��z��������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h0nj h�   hh�j�g������u̃}� u1�����    j h�   hh�h8�h0n�bz��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj ��y�����Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj �y�����E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPhx��kp�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhx��	p�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�j h  hh�j�td������u̃}� u1�~���    j h  hh�h4�h��Ow���������  �} t�} v	�E�   ��E�    �U�U�}� u!h��j h  hh�j��c������u̃}� u1�}���    j h  hh�h4�h����v��������j  �MQ�UR�EP�MQ�URh?��n�����E��}� }X3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���M�U���Rh�   �E��P��c�����}��uu3�t	�E�   ��E�    �U�U��}� u!h\�j h  hh�j��b������u̃}� u.�|��� "   j h  hh�h4�h\���u��������m�}� |d�}�t^�}���tU�M���;MsJ�U����E+�9�As��A�M���U����E+E��M���Qh�   �U��E�LPQ��b�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�$j����]���������������̋�U���,�E������E�    3��} ���E�}� u!h�j h9  hh�j�=a������u̃}� u1��z���    j h9  hh�hX�h��t��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!h��j h?  hh�j�`������u̃}� u1�5z���    j h?  hh�hX�h���s��������  �M;M��   ��y����U��EP�MQ�UR�E��P�MQh?��Ok�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9�As��A�U���E���M+ȉM�U���Rh�   �E�M�TAR�k`�����Yy���8"u
�Oy���M�������  �c�;y����U��EP�MQ�UR�EP�MQh?��j�����E�3ҋE�Mf�TA��}��u"�}�u��x���8"u
��x���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9�As
��A�E��	�M���M��U���Rh�   �E��P�_�����}��ux3�t	�E�   ��E�    �U܉U�}� u!h\�j hf  hh�j�^������u̃}� u1�)x��� "   j hf  hh�hX�h\��sq��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9�As��A�M���U����E+E؋M���Qh�   �U��E�LPQ�^�����}� }	�E�������U��UԋEԋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�h����]�����������̋�U����EPj �MQ�UR�EPhն�g�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhն�Ig�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uh�Nj jfh��j�N[������u̃}� u0��t���    j jfh��h��h�N�,n�����   �  3�;U��؉E�uh��j jgh��j��Z������u̃}� u0�}t���    j jgh��h��h����m�����   �  3ҋEf��}�tK�}���tB�}v<�M��9�As��A�U��	�E���EԋM���Qh�   �U��R�[����3��} ����;E��ىM�uhP�j jih��j�'Z������u̃}� u0�s��� "   j jih��h��hP��m�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uh�j jjh��j�Y������u̃}� u0�<s���    j jjh��h��h��l�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!h��j h�   h��j�X������u̃}� u0�)r��� "   j h�   h��h��h���sk�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�e�����]�����������������̋�U��j �EP�MQ�UR�EP�4���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!h�Nj h>  h��j�V������u̃}� u3�o���    j h>  h��h��h�N��h�����   �A  3�;U���؉E�u!h��j h?  h��j�U������u̃}� u3�.o���    j h?  h��h��h���xh�����   ��  3ҋE�f��}��tK�}����tB�}�v<�MЃ�9�As��A�U��	�EЃ��E̋M���Qh�   �Uԃ�R�U����3��} ����;E���ىM�u!hP�j hA  h��j��T������u̃}� u3�cn��� "   j hA  h��h��hP��g�����"   �  �}r�}$w	�E�   ��E�    �EȉE܃}� u!h�j hB  h��j�PT������u̃}� u3��m���    j hB  h��h��h��+g�����   �  �E�    �UԉU��} t0�-   �M�f��U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ�m���E�U3�PR�MQ�UR�l���E�U�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} w�} v�M�;M�r��U�;U�rn3��M�f��U�;U���؉E�u!h��j hf  h��j�S������u̃}� u0�l��� "   j hf  h��h��h����e�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�"���]����������������̋�U����  ��A3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���[���E�    �j���E�3Ƀ} �������������� u!h��j h  h�j�P������u̃����� uF�Gj���    j h  h�h��h���c����ǅ<��������M���j����<����  3��} �������������� u!hoj h  h�j�1P������u̃����� uF�i���    j h  h�h��ho�	c����ǅ8��������M��=j����8����!  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U����  ������ ��  �������� |%��������x��������x�����,����
ǅ,���    ��,�����������������������И�����������������(�����(����*  ��(����$�Dg	�E�   ������Q�UR������P�h  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ��������$�����$����� ��$�����$���wL��$�����|g	�$�dg	�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�pe�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�e�����Ẽ}� }�E�������M�k�
�������DЉE��  �������� ����� �����I�� ����� ���.�  �� ������g	�$��g	�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  �������h	�$��g	�M���0  u	�U��� �U��E�   �EP�Mc����f�������M��� tW���������   ������ƅ���� �M��K��P�M��K��� ���   Q������R������P�c������}�E�   �f������f�������������U��E�   �  �EP�b���������������� t�������y u��N�U��E�P�N�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ����������������MQ��a�����E��U��� ��   �}� u��N�E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M��I��P�������Q�K������t������������������������������d�}� u	��N�M��E�   �U���|�������������������������t��|������t��|�������|����ɋ�|���+U����U��  �EP��`������x�����V������   3�tǅ���   �
ǅ���    �������t�����t��� u!h@�j h�  h�j�$I������u̃�t��� uF�b���    j h�  h�h��h@���[����ǅ4��������M��0c����4����  ��  �M��� t��x���f������f����x�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h�j�Ḿ�]  Q�BA�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��G��P�U�R�E�P������Q�U�R�E�P��h���Q��AR�ܑ�Ѓ��E�%�   t%�}� u�M���F��P�M�Q��AR�ܑ�Ѓ���������gu)�M���   u�M��F��P�U�R��AP�ܑ�Ѓ��M����-u�E�   �E��M����M��U�R�oJ�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�M������X�����\����   �U���   t�EP�]M������X�����\����   �M��� tB�U���@t�EP�a]��������X�����\�����MQ�E]���������X�����\����=�U���@t�EP�]�������X�����\�����MQ�]����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R�k^����0��d����E��RP��T���P��P���Q��\����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �]  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��B��P�M��B������   R��H���P������Q�Z������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��L���Rj �  ���}� tj�E�P�TQ�����E�    �"�����������0����M��\����0����M�3��;����]Ð�Y	 Z	SZ	�Z	[	"[	e[	�\	�Z	�Z	�Z	�Z	�Z	�Z	 �I �[	�\	�[	�\	�\	 �Z`	�\	#^	 b	�]	r`	�\	�a	c_	gb	b	6^	b	,b	e	   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�O�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U���@�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!hoj h�   hh�j�g:������u̃}� u1��S���    j h�   hh�h��ho�BM��������V  3Ƀ} ���MЃ}� u!hx�j h�   hh�j��9������u̃}� u1�S���    j h�   hh�h��hx���L���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P�T�����E��} u�E��   �M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �L�����EȋE��H���MċU��EĉB�}� |!�M��� 3�%�   �E��M�����E����M�Qj �DL�����E��E���]��������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�oN����]�������������������̋�U��EP�MQ�UR�EP�=N����]�����������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!hoj h�  hh�j�7������u̃}� u.�(Q���    j h�  hh�h��ho�rJ��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQhx���H����]������������������̋�U��EP�MQ�URhx��H����]����������������̋�U��EPj �MQhն�aH����]������������������̋�U��EP�MQ�URhն�/H����]����������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]������������������̋�U����E��t
�-�R�]���M��t����-�R�]������U��t
�-�R�]���E��t	�������؛�M�� t���]����]�������������������������̋�U��Q�=�� t�]���E�    �E���]�������������̋�U��j�hp2h�d�    P���SVW��A1E�3�P�E�d�    �e�=�� ��   �E��@tp�=�R tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe���R    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]�������������������������������������������������������̋�U��Q�=�� t�]��e���U���]�����������������̋�U��Q�=�� t�4���E��E���?�E���E�    �E���]����������������̋�U��Q�=�� t�X4���E��E���?�E���?����E�    �E���]���������������������������̋�U����=�� t8�4���E��E#E�M��#M���E��U������U��U��E�P�1������E�    �E���]�������������������������̋�U��Q�3���E��E��?E��E��M�Q�J1������]����������������������̋�U���@��A3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �M�y ��  �U�z u+�E��Ph  �M�Q0Rj �E�P�G6������t�"  j^h��jj�+�����E�jbh��jjh�  �J�����E�jdh��jjh�  �J�����E�jfh��jjh�  �fJ�����E�jhh��jjh  �KJ�����E�}� t�}� t�}� t�}� t�}� u�}  �M��    �U�U��E�    �	�E����E��}�   }�M��U���E����E��ۍM�Q�U�BP�����u�&  �}�v�  �M܉Mă}�~S�U�U��	�E����E��M����t8�E��H��t-�U���E��	�M����M��U��B9E��M�M�� ���j j �U�BP�Ḿ�   Qh   �U�Rjj ��=���� ��u�  j �E�HQh�   �Uȁ   Rh�   �E��Ph   �M�QRj �>����$��u�E  j �E�HQh�   �U��   Rh�   �E��Ph   �M�QRj �@>����$��u�  3��M�f���   �U��B �E��@ �M�Ɓ�    �U�Ƃ�    �}�~]�E�E��	�M����M��U����tB�M��Q��t7�E���M��	�U����U��E��H9M�� �  �E��M�f��A   ���h�   �Ú�   R�E�P�9����j�Mȁ�   Q�U�R�h9����j�E�   P�M�Q�Q9�����U���    ��   �E���   Q�(�����   3�uj j h�   hX�j�.������u�j�M���   ���   R�>����j�E���   ��   Q��=����j�U���   -�   P��=����j�M���   R�=�����E��    �M�UЉ��   �E�   �M���   �Ú��   �E���   �Mȁ��   �U���   �E��   �M���   �U�Eĉ��   j�M�Q�E=����3���   j�U�R�0=����j�E�P�"=����j�M�Q�=����j�U�R�=����j�E�P��<�����   �   �   �M���    tA�U���   P�(���u-�M���    w!h�j h�   hX�j�/-������u̋Eǀ�       �Mǁ�       �0��E���   ����U���   �8��M���   �Uǂ�      3��M�3���&����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����d4���E��E��Hl�M��U�;LKt�E��Hp#�Hu�Q;���E��U����   ��]�������������������������̋�U��Q�} u
��A���E���E����   �U��E���]���������������������̋�U�����3���E��E��Hl�M��U�;LKt�E��Hp#�Hu�:���E��U��B��]����������������������������̋�U����d3���E��E��Hl�M��U�;LKt�E��Hp#�Hu�Q:���E��U��B��]����������������������������̋�U����3���E��E��Hl�M��U�;LKt�E��Hp#�Hu��9���E��E�����]����������������������������̋�U��3�]��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^���������������������������̋�U��Q�E�    �} u3��S  �}��   �	�E����E��M��9M���   �U���U�E���E�M�Q���t�E�H��U�B�;�t�M�A��U�J�+���   �U�B���t�M�Q��E�H�;�t�U�B��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��X�����	�E����E��M�;Ms>�U���t�M��E�;�t�U��M�+���E���E�M���M�3���]������������������������������������������������������������������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U���(�E�E��M�M��U�U��}��g  �E��$���	�M�Q�U�R��  ���E�}� t�E�E��s�M���Q�U���R��  ���E�}� t�E�E��F�M���Q�U���R�  ���E�}� t�E�E���M���Q�U���R�  ���E�E�E�M�M�E���   �U�R�E�P�Y  ���E�}� t�M�M��F�U���R�E���P�2  ���E�}� t�M�M���U���R�E���P�  ���E܋M܉M��E��i�U�R�E�P��   ���E�}� t�M�M���U���R�E���P��   ���E؋E��*�M�Q�U�R�   ���3���EP�M�Q�U�R�  ����]Ðw�	e�	&�	��	�	�����������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��+�P�   ����]�����������������̋�U��} t3��} ���D ��E�E]����������������̋�U����} �R  �EP�MQ�Q	  ���E��}� t�E��O  �U��R�E��P�*	  ���E��}� t�E��(  �M��Q�U��R�	  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�g  ���E��}� t�E��e  �U��R�E��P�@  ���E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$��	�U��R�E��P��  ���E��}� t�E���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��}  �U��R�E��P�X  ���E��}� t�E��V  �M��Q�U��R�1  ���E��}� t�E��/  �E��P�M��Q�
  ���E��}� t�E��  �U��R�E��P��  ���E��}� t�E���  3���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��  �U��R�E��P�g  ���E��}� t�E��e  �M��Q�U��R�@  ���E��}� t�E��>  �E��P�M��Q�  ���E��}� t�E��  �U��	R�E��	P��  ���E��}� t�E���  �M��Q�U��R��  ���E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�b  ���E��}� t�E��`  �E��P�M��Q�;  ���E��}� t�E��9  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���E��}� t�E���  �E��
P�M��
Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���  �E��P�M��Q�]  ���E��}� t�E��[  �U��R�E��P�6  ���E��}� t�E��4  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���   �U��R�E��P��  ���E��}� t�E��   �M��Q�U��R�  ���E��}� t�E��   �E��P�M��Q�s  ���E��}� t�E��t�U��R�E��P�o������E��}� t�M��M��F�U��R�E��P�H������E��}� t�M��M���U��R�E��P�!������E��M��M�E��3���]Ë�1�	I�	u�	��	
�	"�	N�	z�	�	��	'�	S�	��	ԇ	 �	,�	��	��	و	�	n�	��	��	މ	G�	_�	��	��	 �	8�	d�	��	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��;�tK�E�E��M�M�U�R�E�P�������E�}� t�M�M���U���R�E��P�\������E�E��3���]�������������������������������������������̋�U��� �E�E��M�M��U��E��
;��   �U�U��E�E�M�Q�U�R��������E�}� t�E�E��s�M���Q�U��R�������E�}� t�E�E��F�M���Q�U��R�������E�}� t�E�E���M���Q�U��R�n������E��E��E�M�M�E��3���]�����������������������������������������������������������������̋�U�����"���   �E��} u�E�P�\  ���  �M��U��E��@�M��A�U��z t#�E��H���t�E���PjhP���  ���M��A    �U��: ��   �E�������   �E��x t�M��Q���t�M�Q�O  ����U�R�	  ���E��x uG�M�Qj@h���u  ����t0�U��z t�E��H���t�E�P��  ����M�Q�1	  ���0�U��z t�E��H���t�E�P�  ����M�Q�?  ���U��z u3��N  �} t�E�   �E���E�    �M�Q�U�R�U  ���E��}� t!�}���  t�}���  t�E�P�����u3���   j�M��QR� ���u3���   �} t&�E�M�f�Qf��E�M�f�Qf�P�Ef�M�f�H�} ��   �U�=  u4j h1  h�h|h` hD j@�MQ�2����P�U#����� j@�URh  �E��HQ�����u3��Bj@�U��@Rh  �E��HQ�����u3��j
j�U�   R�E�P��+�����   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�;Eb�}� t\�E�E�+����E��M��U��P�M�R�/�����E�}� u�E��M�T��E���}� }�M����M�	�U����U��3��}� ����]�����������������������������������̋�U��Q�E�Q�A����3҃��E�P�M�QR�$����3Ƀ����U�J�E�@    �M�y t	�E�   ��U�P��  ���E��M�U��Qjh �	���E�H��   t�U�B%   t�M�Q��u
�E�@    ��]����������������������������������������������������������̋�U���   ��A3ŉE������   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �  �E�P��|����QR��-�������r  jx�E�P��|����Q��ҁ������  R��x���P�����u��|����A    �   �G  �U�R��|����Q�a-������u:��|����B  ��|����A��|�����x����B��|�����x����Q��   ��|����H����   ��|����z tt��|����HQ�U�R��|����Q�O#������uQ��|����B����|����A��|�����x����B��|����R�������|���;Au��|�����x����B�E��|����Q��u7��x���P��  ����t$��|����Q����|����P��|�����x����Q��|����H��   ��   ��  jx�U�R��|����H��Ɂ������  Q��x���R�����u��|����@    �   �  �M�Q��|����P��+�������
  ��|����Q��   ��|����P��|����y t7��|����B   ��|����A��|����z u��|�����x����H�   ��|����z tl��|����Q�`������|���;BuP��|���Pj��x���Q��  ����t2��|����B   ��|����A��|����z u��|�����x����H�2��|����B   ��|����A��|����z u��|�����x����H�   ��|����z ut��|����x th�M�Q��|����P�*������uO��|���Qj ��x���R�C  ����t3��|����H��   ��|����J��|����x u��|�����x����Q��|����@��������M�3��
����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�Q�����3҃��E�P�M�y t	�E�   ��U�P��  ���E��M�U��Qjh�	���E�H��u
�U�B    ��]��������������������������������������������̋�U���   ��A3ŉE�����   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �  �E�P��|����R��'������u`��|����x u��|���Qj��x���R�y  ����t3��|�����x����H��|�����x����B��|����Q����|����P�   ��|����y ut��|����z th�E�P��|����R�F'������uO��|���Pj ��x���Q��  ����t3��|�����x����B��|�����x����Q��|����H����|����J��|����@��������M�3��p����]� ������������������������������������������������������������������������������������������������������̋�U��E�HQ�a����3҃��E�PjhP�	���M�Q��u
�E�@    ]��������������������������̋�U���   ��A3ŉE�����   ��|����EP�B  ����x���jx�M�Q��|����B���%���  P��x���Q�����u��|����B    �   �s�E�P��|����QR�y%������uF��x���P��  ����t3��|�����x����Q��|�����x����H��|����B����|����A��|����B��������M�3������]� ������������������������������������������������������������������̋�U��Q�E�H��  �U�J���E��E�M��H�U�E��B��]�������������������������̋�U��Q�} t�E���th4�UR�������u0j�E�Ph  �M�QR�����u3��Y�}� u����K�Fh0�EP�K������u"j�M�Qh   �U�BP�����u3����MQ�#�����E��E���]��������������������������������������������������������̋�U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E, ;�u3���ظ   ��]����������������������̋�U���V�E%�  �ȁ�   �щU�j�E�Ph   �M�Q�����u3��9�U;U�t,�} t&�E�Q��   �����U�P������;�u3���   ^��]������������������������������������̋�U����E�    �E��M��U��E���E��tM�M���a|�U���f�E���'�E���M���A|�U���F
�E����E��M����U��DЉE�뚋E���]������������������������������������̋�U����E�    �E��M��U���U�E���A|	�M���Z~�U���a|%�E���z�M����M��U��E��M���M���E���]�������������������������̋�U���EP�MQ�u����]�������̋�U��Q�E=��  u3��G�M��   }�U�<O�P�M#��&�U�Rj�EPj����u3�f�M��E��U#�]��������������������������������̋�U���EP�MQ������]�������̋�U����d����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR��	�����   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�i   �� �   ��]���������������������������������������������������������������������������������������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}������E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  ������    u��  ������   �E�������   �M�E�j�UR�������t��M���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u���������    ty�t�����   �E��f��ǀ�       �M�Q�UR��  ������t�C�M�Q�  ���Ѕ�t+j�EP������h<�M�����h�2�M�Q��������U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP������E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q��������u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�  ��,�	���D���������M��tj�UR�<�����E�����   �M��������!���   �E�x ��   �M�QR�EP��  ���ȅ���   ������   �U�������   �E���
���M���   ��
���U���   �}$ u�EP�MQ������UR�E$P����j��MQ�UR�EP������M�QR�C  ���
���M���   �
���U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP�  �� ������>
�����    u�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M��EP�M��_���M��P�E���]� ��������̋�U��Q�M��E�� P�M������]������������������̋�U��Q�M��M�����E��t�M�Q������E���]� �����������������̋�U��Q�M��EP�M��M���M��P�E���]� ��������̋�U���V�E�8  �u�c  ������    tW������`��9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�f������t��   �M�y t��#����U�R�E�P�MQ�U R�EP�}�����E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������������������������������������������������������������������������������������������������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�v ������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����������������������������������������������������̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@�'��ǀ�       ����������    ~����   �E�M����E�3��3���]�������������������������������������̋�U��j�h�2h�d�    P���SVW��A1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E��X���   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}������M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R�����E�    ��E�P������Ëe��E�    �M��M��f����E������   �)������    ~����   �EԋUԋ���MԉËU�;Uu�������E�M�H�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����E�E��}  t�M Q�UR�E�P�MQ������}, u�UR�EP�����MQ�U,R����E$�Q�UR�EP�M�Q�������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�T   ���E��}� t�EP�M�Q�p�����]�������������������������������������������������������̋�U��j�h(3h�d�    P���SVW��A1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R��������E�������   �E��}�����   �M��o���U���   �a���M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP������E��E�    ��   �M�Q�N  ��Ëe����ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�M������E�    �E�    �E������E�    �   �   �M�U��Q��E�P�����������Mȉ��   ������Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP�	������t�M�Q�UR�O����ËEЋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u�m���ǀ     �   ��3���]�����������������������������������̋�U��j�hX3h�d�    P���SVW��A1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR�^�������t9j�E�P��������t'�M��U�B��M��Q�U��P�J������M��������@  �U���txj�M�QR���������tYj�E�P�-�������tG�M�QR�E�HQ�U�R�������E�xu"�M��9 t�U��R�E��Q��������U����7����   �E�x uZj�M�QR�{�������t>j�E�P��������t,�M�QR�E��P�M�QR�j�����P�E�P��������������[j�M�QR�!�������tAj�E�P�R�������t/�M�QR��������t�E���t	�E�   ��E�   ��t����E�������   Ëe��\����E������E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hx3h�d�    P���SVW��A1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�<�����E��}�t�}�t+�R�U��R�E�HQ������P�U�BP�M�Q������)j�U��R�E�HQ�[�����P�U�BP�M�Q�����E�������   Ëe������E������M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h�3h�d�    P��SVW��A1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR�����E�������E�����Ëe������E������M�d�    Y_^[��]�������������������������������������������������̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]������������������������̋�U������3Ƀ��    ����]������̋�U���(�} u3���  �E��M��} t�U�B����   �M��9MOC�t�U��:RCC�t�E��@uz�M��9csm�uK�U��zuB�E��x �t�M��y!�t�U��z"�u�E��x u��������    u3��I  ������   �E܋M܋���E܉�   �%  �M��9csm��  �U��z�  �E��x �t�M��y!�t�U��z"���   �E��x u#�U������    u3���   �@������   �M��U�U�E�E��M���   ��M��U��B�H���M�U��B�H��U���E����E��M���M�}� ~d�U��E��M��QR�E�P�M�Q��������t?������   �E؋U؋���M؉�} t�U�R�E�P�MQ�U�R������   ��3���]�����������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E��M����M�U���U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u�v������   �E��M��QR�E�P�������E��R����M􋐈   ��B����M����   ��2����M����   ��U�������E�� ���������   �E�M����E���������    }�����ǀ�       �   ��]������������������������������������������������������������������������������������̋�U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!�!����   �E��U�����M���   �3���]����������������������������������������������̋�U����E�E��M����M�U���U��E�8��G  �M�Q�������} ��   �������   �:csm�u~�w������   �xum�f������   �y �t(�R������   �z!�t�>������   �x"�u1�*������   �QR��������tj�������   P���������������   �9csm�um��������   �zu\��������   �x �t(��������   �y!�t�������   �z"�u �} t�����   �E��E�����U��
�y����M����   �i����M�����   ��]���������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U��j�h�3h�d�    P��SVW��A1E�3�P�E�d�    �e��E�    �M�U�E�������E�P������Ëe��E������M�d�    Y_^[��]��������������������������������������������̋�U��j�h�3h�d�    P��SVW��A1E�3�P�E�d�    �e��E�    �EP�U���E�������M�Q�������Ëe��E������M�d�    Y_^[��]����������������������������������������̋�U��j�h�3h�d�    P��SVW��A1E�3�P�E�d�    �e��E�    �EP�U�E�������M�Q�`�����Ëe��E������M�d�    Y_^[��]�������������������������������������������̋�U��j�h4h�d�    P��SVW��A1E�3�P�E�d�    �e��E�    �EP�MQ�UR�EP�U�E�������M�Q������Ëe��E������M�d�    Y_^[��]�����������������������������������������������̋�U����} t������} u�����E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR��������t�E���뀊E��]������������������������������������������������������������̋�U��j�h��
d�    PQSVW��A3�P�E�d�    �e��1������    u������E�    �A����$�����M���   j j �~����E������)�	��E������b����M�d�    Y_^[��]������������������������������������������������̋�U��Q�E�    �	�E����E��M�U�;}'h�R�E����M�Q�L��������t����2���]���������������������������������̋�U����} t������E��M�}� t������U�:csm�u/�E�xu&�M�y �t�U�z!�t�E�x"�u��H����M�Q�B���E��M�Q�B��M���U����U��E����E��}� ~0�M���U��E��H��Q�M����P���������u�   ��3���]�����������������������������������������������������������U���SQ�E���E��EU�u�M�m��}���VW��_^��]�MU���   u�   Q�[���]Y[�� �������������������̋�U�����A3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ��������UR��������E�P�MQ�������UR��������E��M��E�    �E�    �U�R�EP��������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR�E�����f�E�f��f�E��؋Mf�U�f�Q
�M�3��U�����]����������������������������������������������������������������������������������������������̋�U��=�m uj �EP�MQ�URhPK�:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h�
d�    P��H��A3�P�E�d�    �EP�M��@����E�    �} t�M�U�3��} ���Ẽ}� uhLj j^h�j��������u̃}� uD�����    j j^h�h�hL��������E�    �E������M��,����E��  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uh`j j_h�j��������u̃}� uD�����    j j_h�h�h`�f������E�    �E������M������E��v  �M�M��E�    �U���E�M����M��M��t�����t0�M��h�������   ~�M��U���Pj�E�P�������E��j�M�Q�M��1���P��������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} |�}t�}$~.�} t�U�E��E�    �E������M������E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M����M��U���E�M����M�����3��u�E�j�U�R�M�����P�f�������t�E��0�E��Qh  �M�Q�M�����P�;�������t0�U��a|�E��z�M�� �M���U�U��E���7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M���U�E����E��!����M����M��U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4������ "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U���E��t�M��ىMЋUЉU��E������M������E��M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U��=�m uj�EP�MQ�URhPK��������j�EP�MQ�URj �n�����]�������������������������̋�U��j�EP�MQ�UR�EP�4�����]���������������̋�U��=�m uj �EP�MQ�URhPK�:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h8�
d�    P��lVW��A3�P�E�d�    �EP�M�������E�    �} t�M�U�3��} ���E��}� uhLj j^h�j���������u̃}� uN�m����    j j^h�hlhL�������E�    �E�    �E������M�������E��U��<  �} t�}|�}$~	�E�    ��E�   �U��U��}� uh`j j_h�j�<�������u̃}� uN������    j j_h�hlh`�������E�    �E�    �E������M��C����E��U��  �M�M��E�    �E�    �U���E�M����M��M�������t0�M���������   ~�M������Pj�E�P�&������E��j�M�Q�M������P�������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E����E��M���U�E����E��E�RPj�j�������E�U�j�M�Q�M������P��������t�U��0�U��Th  �E�P�M�����P�T�������t0�M��a|�U��z�E�� �E���M�M��U���7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u^�U�;U�uV�u�3��E�RPj�j������u��}��E��U��E�;E�w.r�M�;M�w$�E�RP�U�R�E�P�����M�3��։EĉU���U���U�} u��E���M�U����U�������E����E��M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�v���� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M���U��t�E��؋Mȃ� �ىEĉMȋUĉU��EȉE��E������M������E��U��M�d�    Y_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�t�����]���������������̋�U��=�m uj�EP�MQ�URhPK�:�������j�EP�MQ�URj ������]�������������������������̋�U��j�EP�MQ�UR�EP�������]���������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����'  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tE�U�;U�u.�E�H��  ����ًU��  �����;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���(  ��A3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T�������ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �������|���3Ƀ} ����0�����0��� u!h��j h  h�j��������u̃�0��� uI�����    j h  h�h(h���������ǅ ���������T��������� �����7  �E��,�����,����Q��@��   ��,���P��������(�����(����t-��(����t$��(�������(������������\����
ǅ\���B��\����H$�����х�uV��(����t-��(����t$��(�������(������������X����
ǅX���B��X����B$�� ���ȅ�tǅT���    �
ǅT���   ��T�����$�����$��� u!h��j h  h�j��������u̃�$��� uI�����    j h  h�h(h���d�����ǅ����������T��������������T6  3Ƀ} ���� ����� ��� u!hoj h  h�j��������u̃� ��� uI�����    j h  h�h(ho�������ǅ����������T����
�����������5  ǅL���    �E������ǅ@���    ���@�������@�����@����q5  ��@���u������ u�Z5  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Uǅ��������ǅ��������ǅp�������ǅ���������E���G�����G����E���E����1  ��L��� ��1  ��G����� |%��G�����x��G�����(����P����
ǅP���    ��P�����H�����H���k�	��8�����H����8�����8�����  �E���%��  �������u\j
��t���R�EP��������~9��t������$u+��@��� uh@  j ������P������ǅ����   �
ǅ����    �������)  j
��t���Q�UR�R���������������t������E��@��� ��   ������ |#��t������$u������d}ǅL���   �
ǅL���    ��L������������� u!hxj hQ  h�j��������u̃���� uI�����    j hQ  h�h(hx�������ǅ����������T����'�����������2  ������;�x���~��������H������x�����H�����H�����x����   ��8�����   3�tǅD���   �
ǅD���    ��D������������� u!h j h]  h�j�6�������u̃���� uI������    j h]  h�h(h ������ǅ����������T����?�����������1  ��8�����@�����@�����.  ��@����$� 
��@��� u	������t��@���u�������u�.  ǅ����    ��T��������P��G���R�����������   ��L���P�MQ��G���R�9A  ���E���G����U���U��G�������؉����u!h��j h�  h�j��������u̃���� uI�����    j h�  h�h(h���������ǅ����������T���������������0  ��L���R�EP��G���Q�@  ���-  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �P-  ��G�����<�����<����� ��<�����<���wi��<�����X
�$�@
���������������D���������������3���������������"�������   ����������������������,  ��G�����*��  ������ u�EP��������������^  j
��t���Q�UR����������������t������E��@��� ��  ������ |#��t������$u������d}ǅ8���   �
ǅ8���    ��8������������� u!hhj h�  h�j���������u̃���� uI�g����    j h�  h�h(hh������ǅ����������T���������������.  ������;�x���~��������4������x�����4�����4�����x����������������� uE��������Ǆ����   ����������G������������������������������   ������P��G���Qj��������������P����������؉����u!h�
j h�  h�j��������u̃���� uI�0����    j h�  h�h(h�
�z�����ǅ����������T��������������j-  �\*  �+������������������������Q������������������ }���������������������؉������������k�
��G����DЉ�������)  ǅd���    ��)  ��G�����*��  ������ u�UR���������d����^  j
��t���P�MQ�)���������p�����t������U��@��� ��  ��p��� |#��t������$u������d}ǅ0���   �
ǅ0���    ��0������������� u!h
j h�  h�j���������u̃���� uI�����    j h�  h�h(h
�������ǅ����������T���������������+  ��p���;�x���~��p�����,������x�����,�����,�����x�����p����������� uE��p�����Ǆ����   ��p�������G�����������p������������������   ������R��G���Pj��p�����������R�����������؉� ���u!h`	j h�  h�j��������u̃� ��� uI�L����    j h�  h�h(h`	������ǅ����������T���������������*  �x'  �+��p�����������������������P��������d�����d��� }
ǅd����������d���k�
��G����DЉ�d����'  ��G�����(�����(�����I��(�����(���.�B  ��(������
�$�l
�U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅ8���    �*����"�������� �������������   �������%  ��G�����$�����$�����A��$�����$���7��"  ��$������
�$��
��������0  u������   ��������������  �_  ǅ����    ������ u�UR�=�����f��<�����  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!h 	j h�  h�j蟽������u̃����� uI�-����    j h�  h�h(h 	�w�����ǅ����������T��������������g'  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�����u!hXj h�  h�j菼������u̃����� uI�����    j h�  h�h(hX�g�����ǅ����������T��������������W&  �   �,��������������������������P�E�����f��<�����<���Qh   ��P���R������P������������������ t
ǅl���   �*  ������ u�MQ������f��������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h 	j h�  h�j�J�������u̃����� uI������    j h�  h�h(h 	�"�����ǅ����������T����S����������%  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�F���������؉�����u!h�j h�  h�j�:�������u̃����� uI������    j h�  h�h(h�������ǅ����������T����C����������$  �j  �,��������������������������R������f��������������P���ǅ����   ��P����������  ������ u�UR���������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h 	j h�  h�j��������u̃����� uI�����    j h�  h�h(h 	�������ǅ����������T���������������"  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�����u!hj h�  h�j� �������u̃����� uI�����    j h�  h�h(h�������ǅ����������T����	�����������!  �0  �+��������������������������P������������������� t�������y u#��N������������P軺�����������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������a  ������%0  u��������   ��������d����uǅ���������d������������������������� u�MQ���������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h 	j h6  h�j��������u̃����� uI�����    j h6  h�h(h 	�������ǅ����������T���������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�����u!hj h:  h�j� �������u̃����� uI�����    j h:  h�h(h�������ǅ����������T����	�����������  �0  �+��������������������������R�������������������%  tx������ u��N������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������i������ u��N����������������������������������������t���������t���������������ɋ�����+������������  ������ u�UR���������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h 	j h�  h�j��������u̃����� uI�����    j h�  h�h(h 	�������ǅ����������T���������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�����u!hj h�  h�j���������u̃����� uI�����    j h�  h�h(h�������ǅ����������T���������������  �+  �+��������������������������P��������������ž������   3�tǅ���   �
ǅ���    ����������������� u!h@�j h�  h�j��������u̃����� uI�����    j h�  h�h(h@��������ǅ����������T����#�����������  �J  �������� t������f��L���f����������L����ǅl���   �  ǅh���   ��G����� ��G�����������@��������������  ��@��� ��  ������ |������d}ǅ���   �
ǅ���    ����������������� u!h 	j h�  h�j��������u̃����� uI�v����    j h�  h�h(h 	�������ǅ����������T���������������  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�����u!hpj h�  h�j��������u̃����� uI�s����    j h�  h�h(hp������ǅ����������T���������������  �  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��G�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Zh�  h�j��d�����]  R�7����������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�U���U�E�H��P��������������  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!h 	j h  h�j�<�������u̃����� uI������    j h  h�h(h 	������ǅ����������T����E����������  ��@���t!h0j h  h�j���������u̋����������������������������������������H��P���������������T����ԫ��P��h���P��d���Q��G���R��P���P������Q������R��AP�ܑ�Ѓ���������   t-��d��� u$��T����u���P������R��AP�ܑ�Ѓ���G�����gu3��������   u%��T����7���P������P��AQ�ܑ�Ѓ����������-u!��������   ��������������������������P��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ��������   t ƅ����0��4�����Q������ǅ����   �*ǅ����   ��������   t��������   ������������% �  �#  ������ u�MQ�˱������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u!h 	j h�  h�j�2�������u̃�l��� uI������    j h�  h�h(h 	�
�����ǅ����������T����;�����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�.���������؉�h���u!h�j h�  h�j�"�������u̃�h��� uI�����    j h�  h�h(h��������ǅ����������T����+�����������  �R  �1����������������d�����d���R�ί������x�����|�����
  ������%   �#  ������ u�MQ藯������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������`�����`��� u!h 	j h�  h�j���������u̃�`��� uI�����    j h�  h�h(h 	�ֺ����ǅ����������T���������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�����������؉�\���u!h�j h�  h�j��������u̃�\��� uI�|����    j h�  h�h(h��ƹ����ǅ����������T���������������  �  �1����������������X�����X���R蚭������x�����|�����  �������� �a  ��������@�'  ������ u�UR臽��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������T�����T��� u!h 	j h�  h�j軥������u̃�T��� uI�I����    j h�  h�h(h 	蓸����ǅ����������T����Ŀ���������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R跭��������؉�P���u!h�j h�  h�j諤������u̃�P��� uI�9����    j h�  h�h(h�胷����ǅ����������T���贾���������s  ��  �3����������������L�����L���P舻��������x�����|����&  ������ u!�MQ�`����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������H�����H��� u!h 	j h�  h�j蒣������u̃�H��� uI� ����    j h�  h�h(h 	�j�����ǅ����������T���蛽���������Z  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q莫��������؉�D���u!h�j h�  h�j肢������u̃�D��� uI�����    j h�  h�h(h��Z�����ǅ����������T���苼���������J  �  �5����������������@�����@���R�_����������x�����|����V  ��������@�%  ������ u�MQ�&��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������<�����<��� u!h 	j h  h�j�[�������u̃�<��� uI�����    j h  h�h(h 	�3�����ǅ����������T����d����������#  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�W���������؉�8���u!h�j h  h�j�K�������u̃�8��� uI�ٹ���    j h  h�h(h��#�����ǅ|���������T����T�����|����
  �{  �2����������������4�����4���R�(��������x�����|����"  ������ u�EP������3ɉ�x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������0�����0��� u!h 	j h0  h�j�5�������u̃�0��� uI�ø���    j h0  h�h(h 	������ǅx���������T����>�����x�����  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�1���������؉�,���u!h�j h4  h�j�%�������u̃�,��� uI賷���    j h4  h�h(h��������ǅt���������T����.�����t�����  �U  �3����������������(�����(���R������3ɉ�x�����|�����������@tG��|��� >|	��x��� s3��x����؋�|����� �ى�p�����t�����������   ���������x�����p�����|�����t����������� �  u(������%   u��p�����t����� ��p�����t�����d��� }ǅd���   �%�����������������d���   ~
ǅd���   ��p����t���u
ǅ����    ��O�����������d�����d�������d�������p����t�����   �������RP��t���P��p���Q�1�����0�������������RP��t���R��p���P萴����p�����t���������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�s  ��l��� �B  ��������@t[��������   tƅ����-ǅ����   �:��������tƅ����+ǅ����   ���������tƅ���� ǅ����   ������+�����+�������$�����������u��L���Q�UR��$���Pj �m  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��$���Qj0�  �������� ��   ������ ��   ǅ���    �������� �����������������������������������   �� ���f�f������������Rj�����P�����Q蝴����������� ������� �������� u	����� uǅL��������-��|���P��L���Q�UR�����P�����Q�  ���S����(��|���R��L���P�MQ������R������P�P  ����L��� |'��������t��L���R�EP��$���Qj ��  �������� tj������R�f�����ǅ����    ������8��� t��8���tǅ����    �
ǅ����   ���������������� u!hhj h�  h�j茘������u̃���� uI�����    j h�  h�h(hh�d�����ǅp���������T���蕲����p����T  �������%  ��@��� �  ǅ����    ���������������������;�x�����  �����������������������������������������  �������$�$
���������E�������MQ�������  ���������E�������MQ襨�����_  ���������E�������MQ訮�����;  ���������E�������MQ�S������  ���������E�������MQ�/�������   ���������E�������MQ�<�������   ���������E�������MQ���������h�����l����   3�tǅ����   �
ǅ����    ���������������� u!h�j h.	  h�j�\�������u̃���� uF�����    j h.	  h�h(h��4�����ǅd���������T����e�����d����'������s�����L�����`�����T����<�����`����M�3��ُ����]Ë�8�	f�	��	J�	�	.�	��	`�	�	#�	�	��	6�	E�	 �I i�	9�	-�	J�	[�	 �m�	��	�	��	h�	��	��	~�	m�	�	��	;�	��	��	}
   	
B
f
�
�
�
�
J

�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP��������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U���<  ��A3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��n����E�    �!����E�3Ƀ} �������������� u!h��j h  h�j�I�������u̃����� uF�ל���    j h  h�h�h���!�����ǅ��������M��U���������#  �E�������������Q��@��   ������P�ٌ�����������������t-�������t$����������������������������
ǅ����B�������H$�����х�uV�������t-�������t$����������������������������
ǅ����B�������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h��j h  h�j�ԁ������u̃����� uF�b����    j h  h�h�h��謔����ǅ��������M������������  3Ƀ} �������������� u!hoj h  h�j�L�������u̃����� uF�ښ���    j h  h�h�ho�$�����ǅ��������M��X���������&  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���  ������ �	  �������� |%��������x��������(���������
ǅ����    ������������������k�	��������H����������������   3�tǅ����   �
ǅ����    ������������������ u!h j ha  h�j��������u̃����� uF�n����    j ha  h�h�h 踒����ǅ��������M�����������  ��������������������  �������$�08
�E�    �M��~��P������R輀��������   ������P�MQ������R�u  ���E��������U���U����������؉�|���u!h��j h�  h�j��~������u̃�|��� uF�l����    j h�  h�h�h��趑����ǅ��������M�����������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK��������h8
�$�P8
�E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�
������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ豔�����Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ���������8
�$�|8
�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ���������8
�$��8
�U���0  u�E�   �E��M���  tUǅx���    �UR谌����f������������Ph   ������Q�U�R�%�������x�����x��� t�E�   �&�EP茒����f��t�����t����������E�   �������U��W  �EP�X�������p�����p��� t��p����y u��N�U��E�P�<~�����E��P�M���   t&��p����B�E���p�����+����E��E�   ��E�    ��p����B�E���p�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������h����MQ腑�����E��U���  te�}� u��N�E��E�   �M���d�����h�����h�������h�����t��d������t��d�������d����ɋ�d���+M����M��[�}� u	��N�U��E���l�����h�����h�������h�����t��l������t��l�������l����ɋ�l���+E��E��  �MQ覐������`���蓆������   3�tǅ����   �
ǅ����    ��������\�����\��� u!h@�j h�  h�j��x������u̃�\��� uF�v����    j h�  h�h�h@��������ǅ ��������M�������� �����  ��  �U��� t��`���f������f����`�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h�j�Ú�]  R�q�����E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���P�����T����M���v��P�E�P�M�Q������R�E�P�M�Q��P���R��AP�ܑ�Ѓ��M���   t$�}� u�M��v��P�U�R��AP�ܑ�Ѓ���������gu*�U���   u�M��bv��P�E�P��AQ�ܑ�Ѓ��U����-u�M���   �M��U����U��E�P�2z�����E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�N}������@�����D����   �U���   t�EP�&}������@�����D����   �M��� tB�U���@t�EP�*���������@�����D�����MQ�����������@�����D����=�U���@t�EP���������@�����D�����MQ�͌����3҉�@�����D����E���@t@��D��� 7|	��@��� s,��@����ً�D����� �ډ�8�����<����E�   �E����@�����8�����D�����<����E�% �  u&�M���   u��8�����<����� ��8�����<����}� }	�E�   ��M�����M��}�   ~�E�   ��8����<���u�E�    �E��E��M̋Ũ��U̅���8����<���t{�E��RP��<���Q��8���R�7�����0��L����E��RP��<���P��8���Q虌����8�����<�����L���9~��L����������L����E���L�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅4����M���u������R�EP��4���Qj �K	  ���U�R������P�MQ�U�R�E�P�|	  ���M���t$�U���u������P�MQ��4���Rj0� 	  ���}� ��   �}� ��   ǅ���    �E���0����M܉�,�����,�����,�������,�������   ��0���f�f������������Pj�� ���Q��(���R�6������������0�������0�������� u	��(��� uǅ���������*�M�Q������R�EP��(���Q�� ���R�{  ���V�����E�P������Q�UR�E�P�M�Q�U  �������� |$�U���t������P�MQ��4���Rj ��  ���}� tj�E�P�������E�    ����������� t������tǅ����    �
ǅ����   ���������������� u!hhj h�  h�j�=q������u̃���� uC�ˊ���    j h�  h�h�hh������ǅ���������M��I�����������������������M��-����������M�3���j����]ÍI �)
�*
�*
/+
|+
�+
�+
-
	+
+
�*
�*
!+
*+
 �I 7,
�,
,
�,
-
 ��0
C-
�.
]2
�-
�0
Y-
;2
�/
�2
V2
�.
M2
i2
D5
   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�}�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��j�h�4h�d�    P���SVW��A1E�3�P�E�d�    �E������E�    j�=d������u����C  j�i�����E�    �E�    �	�E���E�}�@��  �M�<��� �#  �U�����E��	�M؃�@�M؋U����   9E���   �M��Q����   �E؃x uaj
�i�����E�   �M؃y u.h�  �U؃�R�D���u	�E�   ��E؋H���U؉J�E�    �   �j
�Fv����Ã}� u+�E؃�P����M��Q��t�E؃�P����4����}� u-�M��A�U�������E����M�U�+�����E��������}��t��   ��   h�   h�jj@j ������E؃}� ��   �E�M؉����<��� �<��	�E؃�@�E؋M������   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃��������D�U�R�b������u�E������������E������   �j��t����ËE܋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} ��   �E;<���   �M���U���������<�um�=X]uB�M�M��}� t�}�t�}�t�(�URj�����EPj�����MQj����U���E���������U�3����E~��� 	   �k���     �����]�����������������������������������������������������������̋�U��Q�} ��   �E;<���   �M���U���������L����   �U���E���������<�th�=X]u<�U�U��}� t�}�t�}�t�"j j����j j����
j j����E���M�������������3����&}��� 	   �j���     �����]������������������������������������������������������������̋�U����}�u�1j���     �|��� 	   ����2  �} |�E;<�s	�E�   ��E�    �M�M��}� u!h��j h;  h0j�b������u̃}� u<�i���     �B|��� 	   j h;  h0hh���u��������   �E���M���������D
������؉E�u!h�j h<  h0j�0b������u̃}� u9�3i���     �{��� 	   j h<  h0hh�� u���������U���E�����������]����������������������������������������������������������������������������������������������̋�U��j�h(5h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP�H��E��}� u�$�P��^��������q  �}�u�M��@�M���}�u
�U���U��JX���E؃}��u�8z���    �g���     ����#  �E�    �EP�M�Q�[�����U���U�E����M؃��������E�D
�M����U؃��������L$�ဋU����E؃��������L$�E����M؃��������D
$$�M����U؃��������D$�E�   �E������   �K�}� u8�U����E؃��������T����E����M؃��������T�M�Q��[����Ã}� t�U؉U���E������EԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hH5h�d�    P���SVW��A1E�3�P�E�d�    �E���M��������M��E�   �U��z u_j
�_�����E�    �E��x u,h�  �M���Q�D���u�E�    �U��B���M��A�E������   �j
��l����Ã}� t!�U���E���������TR����E�M�d�    Y_^[��]��������������������������������������������������������������������������̋�U��E���M���������D
P���]������������������������̋�U��j�hh5h�d�    P���SVW��A1E�3�P�E�d�    j�>^�����E�    �EP�?v����f�E��E������   �j�k�����f�E�M�d�    Y_^[��]���������������������������������������������̋�U��Q�=�V�u��W���=�V�u���  �(j �E�Pj�MQ��VR�����u���  �f�E��]��������������������������������̋�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M��f���M��$[������   t1�M��[��� ���   th j jGh�j�[������u̍M���Z����z u*�} t�Ef��Uf�
�E�   �M��u���E��R  �M��Z��P�E�Q�\��������   �M��Z������   ~R�M��sZ��� �M;��   |=3҃} ��R�EP�M��PZ������   R�EPj	�M��9Z����QR����uB�M��!Z��� �M;��   r�U�B��u"�Dt��� *   �E������M���t���E��   �M���Y������   �U�M���t���E��k�a3��} ��P�MQj�URj	�M��Y��� �HQ����u��s��� *   �E������M��qt���E���E�   �M��]t���E���M��Pt����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�eq����]�������������������̋�U��j�h�5h�d�    P���SVW��A1E�3�P�E�d�    �E�    j�GZ�����E�    �E�   �	�E����E��M�; ���   �Uࡼm�<� t|�M���m���H��   t"�Uࡼm��Q��W�������t	�U���U�}�|=�E���m���� R�P�j�E���m��R��g�����E���m��    �Y����E������   �j�g����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������̋�U��j�h�5h�d�    P���SVW��A1E�3�P�E�d�    �} uj �  ���@�EP�c�����E�    �MQ�,j�����E��E������   ��UR�)i����ËE�M�d�    Y_^[��]������������������������������������������̋�U��} uj �n  ���@�EP�9n������t����+�M�Q�� @  t�EP��`����P�J^��������3�]�����������������������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R�C`����P�U����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����������������������������������������������������̋�U��j�   ��]���������������̋�U��j�h�5h�d�    P���SVW��A1E�3�P�E�d�    �E�    �E�    j�V�����E�    �E�    �	�E����E��M�; ���   �Uࡼm�<� ��   �M���m���H��   ��   �Uࡼm��Q�U�R�M�����E�   �E���m���B%�   te�}u%�M���m��P�`g�������t	�M���M��:�} u4�Uࡼm���Q��t!�E���m��R�"g�������u�E������E�    �   ��E���m��R�E�P�e�����������E������   �j��b����Ã}u�E����E܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������̋�U����} uh`�j j?hXj�JS������u̋M�M��U�R�A]����P��f������u3��  �`���� 9E�u	�E�    ��`����@9E�u	�E�   �3���   ��m����m�M��Q��  t3��   �E��<��m u\j[hjh   ��K�����E�M��U���m�}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U����m�A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]��������������������������������������������������������������������������������������̋�U��Q�} t'�}t!h�j h�   hXj�Q������u̋M�M��} tG�U��B%   t:�M�Q��h�����U��B%�����M��A�U��B    �E��     �M��A    ��]��������������������������������������̋�U��j�h�5h�d�    P���SVW��A1E�3�P�E�d�    �d^���� �E�3��} ���E؃}� uhoj j4h0j�P������u̃}� u+�:j���    j j4h0hho�c��������i�U�R�\�����E�    �E�P��O�����E܋MQ�UR�EP�M�Q�U���E��U�R�E�P�3g�����E������   ��M�Q��a����ËE��M�d�    Y_^[��]�����������������������������������������������������������������������̋�U��EP�MQ�URh���+M����]����������������̋�U��EP�MQ�URh���L����]����������������̋�U��EP�MQ�URhù��L����]����������������̋�U��EPj �MQh���L����]������������������̋�U��EPj �MQh��mL����]������������������̋�U��EPj �MQhù�=L����]������������������̋�U���   ��A3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��Y���E�    ��g���E�3Ƀ} �������������� u!h��j h  h�j��M������u̃����� uF�g���    j h  h�h�h����`����ǅ8��������M��h����8����  3��} �������������� u!hoj h  h�j�qM������u̃����� uF��f���    j h  h�h�ho�I`����ǅ4��������M��}g����4����z  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���h  ������ �[  �������� |%��������x��������(���� ����
ǅ ���    �� ���������������k�	��������H����������������   3�tǅ���   �
ǅ���    ����������������� u!h j ha  h�j�L������u̃����� uF�e���    j ha  h�h�h ��^����ǅ0��������M��f����0����  �����������������*  ������$�\k
�E�   ������Q�UR������P�Y  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ������������������ ����������wL��������k
�$�|k
�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�b�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�a�����Ẽ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  ��������k
�$��k
�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  �������(l
�$��k
�M���0  u	�U��� �U��E�   �EP��_����f�������M��� tW���������   ������ƅ���� �M��G��P�M��G��� ���   Q������R������P�4`������}�E�   �f������f�������������U��E�   �  �EP�I_���������������� t�������y u��N�U��E�P�-K�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ�����������|����MQ�y^�����E��U��� ��   �}� u��N�E��M��������E�    �	�U܃��U܋E�;�|���}L���������t?�M��"F��P�������Q�$H������t������������������������������d�}� u	��N�M��E�   �U���x�����|�����|�������|�����t��x������t��x�������x����ɋ�x���+U����U��  �EP�s]������t����`S������   3�tǅ���   �
ǅ���    �������p�����p��� u!h@�j h�  h�j�E������u̃�p��� uF�C_���    j h�  h�h�h@��X����ǅ,��������M���_����,����  ��  �M��� t��t���f������f����t�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h�j�Ḿ�]  Q��=�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��C��P�U�R�E�P������Q�U�R�E�P��h���Q��AR�ܑ�Ѓ��E�%�   t%�}� u�M��dC��P�M�Q��AR�ܑ�Ѓ���������gu)�M���   u�M��.C��P�U�R��AP�ܑ�Ѓ��M����-u�E�   �E��M����M��U�R� G�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�J������X�����\����   �U���   t�EP��I������X�����\����   �M��� tB�U���@t�EP��Y��������X�����\�����MQ��Y���������X�����\����=�U���@t�EP�Y�������X�����\�����MQ�Y����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R��Z����0��d����E��RP��T���P��P���Q�^Y����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �N  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��>��P�M��>������   R��H���P������Q�1W������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�v  �������� |$�U���t������P�MQ��L���Rj ��  ���}� tj�E�P��M�����E�    �s��������� t������tǅ ���    �
ǅ ���   �� �����<�����<��� u!hhj h�  h�j�>������u̃�<��� uC�W���    j h�  h�h�hh��P����ǅ(��������M��X����(������������$����M���W����$����M�3��7����]�h]
�]
�]
8^
�^
�^
�^
`
^
^
^
�]
*^
3^
 �I A_
�_
_
�_

`
 ��c
L`
�a
�e
�`
�c
``
me
�b
�e
�e
�a
e
�e
�h
   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�UK�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����#  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tA�U�;U�u*�E�H�� ��Ƀ��U�� ��҃�;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ��A3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T�����=��ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    �L����|���3Ƀ} ����0�����0��� u!h��j h  h�j�D2������u̃�0��� uI��K���    j h  h�h�h���E����ǅ,���������T����ML����,����3  3��} ����,�����,��� u!hoj h  h�j�1������u̃�,��� uI�GK���    j h  h�h�ho�D����ǅ(���������T�����K����(����3  ǅL���    �U������ǅ@���    ���@�������@�����@�����2  ��@���u������ u�2  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Mǅ��������ǅ��������ǅp�������ǅ���������Uf�f��D�����D����U���U���K/  ��L��� �>/  ��D����� |%��D�����x��D�����(���������
ǅ����    ��������H�����H���k�	��8�����H����8�����8�����  �U���%��  �������u\j
��t���Q�UR�H4������~9��t������$u+��@��� uh@  j ������R�C0����ǅ����   �
ǅ����    �������)  j
��t���P�MQ��3��������������t������U��@��� ��   ������ |#��t������$u������d}ǅ����   �
ǅ����    ��������(�����(��� u!hxj hQ  h�j��.������u̃�(��� uI�bH���    j hQ  h�h�hx�A����ǅ$���������T�����H����$����40  ������;�x���~���������������x�����������������x����   ��8�����   3�tǅ����   �
ǅ����    ��������$�����$��� u!h j h]  h�j��-������u̃�$��� uI�zG���    j h]  h�h�h ��@����ǅ ���������T�����G���� ����L/  ��8����������������N,  �������$���
��@��� u	������t��@���u�������u�,  ǅ����   ��L���Q�UR��D���P�=  ����+  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �+  ��D����������������� ������������wj���������
�$�ت
���������������E���������������4���������������#�������ʀ   ����������������������	+  ��D�����*��  ������ u�UR�rC�����������`  j
��t���P�MQ�t0��������������t������U��@��� ��  ������ |#��t������$u������d}ǅ|���   �
ǅ|���    ��|����� ����� ��� u!hhj h�  h�j�i+������u̃� ��� uI��D���    j h�  h�h�hh�A>����ǅ���������T����rE���������,  ������;�x���~��������x������x�����x�����x�����x����������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R�'4��������؉����u!h�
j h�  h�j�0*������u̃���� uI�C���    j h�  h�h�h�
�=����ǅ���������T����9D��������+  �(  �+������������������������P�A���������������� }���������������������ډ������������k�
��D����TЉ������2(  ǅd���    �#(  ��D�����*��  ������ u�MQ�@������d����`  j
��t���R�EP�-��������p�����t������M��@��� ��  ��p��� |#��t������$u������d}ǅt���   �
ǅt���    ��t������������� u!h
j h�  h�j�(������u̃���� uI�B���    j h�  h�h�h
�[;����ǅ���������T����B���������)  ��p���;�x���~��p�����p������x�����p�����p�����x�����p����������� uG��p�����Ǆ����   ��p�����f��D���f��������p������������������   ������Q��D���Rj��p�����������Q�A1��������؉����u!h`	j h�  h�j�J'������u̃���� uI��@���    j h�  h�h�h`	�":����ǅ���������T����SA��������(  ��%  �+��p���������������������R�'>������d�����d��� }
ǅd����������d���k�
��D����TЉ�d����_%  ��D�����l�����l�����I��l�����l���.�D  ��l������
�$��
�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������d�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu������   �������ǅ8���    ������#�������� ���������������   ��������#  ��D�����h�����h�����A��h�����h���7�B!  ��h�������
�$�H�
��������0  u�������� ������ǅ����   ������ u�EP�<����f��<�����  ������ |������d}ǅd���   �
ǅd���    ��d������������� u!h 	j hv  h�j�=$������u̃���� uI��=���    j hv  h�h�h 	�7����ǅ���������T����F>��������%  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�"-��������؉����u!h�j hz  h�j�+#������u̃���� uI�<���    j hz  h�h�h��6����ǅ���������T����4=��������$  �  �,���������������� ����� ���Q�:����f��<����������� t_��<���%�   ������ƅ���� ��T�����!��P��T�����!������   R������P��P���Q�V:������}
ǅl���   �f��<���f��P�����P���������ǅ����   �^  ������ u�MQ�Y9������������  ������ |������d}ǅ`���   �
ǅ`���    ��`��������������� u!h 	j h�  h�j�!������u̃����� uI�#;���    j h�  h�h�h 	�m4����ǅ���������T����;���������"  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�z*��������؉�����u!hj h�  h�j� ������u̃����� uI�:���    j h�  h�h�h�[3����ǅ ���������T����:���� �����!  �w  �+��������������������������R�`7���������������� t�������x u#��N������������R�>#�����������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q��������������������  ��������0  u�������� ��������d����uǅ\���������d�����\�����\��������������� u�EP�Z6������������  ������ |������d}ǅX���   �
ǅX���    ��X��������������� u!h 	j h6  h�j�������u̃����� uI�$8���    j h6  h�h�h 	�n1����ǅ����������T����8����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�{'��������؉�����u!hj h:  h�j�������u̃����� uI�7���    j h:  h�h�h�\0����ǅ����������T����7����������  �x  �+��������������������������Q�a4������������������ ��   ������ u��N������������������ǅ����    ���������������������;�����}O���������tB��T�������P�������Q��������t������������������������������v������ u��N������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������'  ������ u�EP�"3������������  ������ |������d}ǅT���   �
ǅT���    ��T��������������� u!h 	j h�  h�j�^������u̃����� uI��4���    j h�  h�h�h 	�6.����ǅ����������T����g5���������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�C$��������؉�����u!hj h�  h�j�L������u̃����� uI��3���    j h�  h�h�h�$-����ǅ����������T����U4���������  �@  �+��������������������������Q�)1�����������'������   3�tǅP���   �
ǅP���    ��P��������������� u!h@�j h�  h�j�k������u̃����� uI��2���    j h�  h�h�h@��C,����ǅ����������T����t3����������  �_  �������� t������f��L���f����������L����ǅl���   �%  ǅh���   ��D����� f��D�����������@��������������  ��@��� ��  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u!h 	j h�  h�j�8������u̃����� uI��1���    j h�  h�h�h 	�+����ǅ����������T����A2���������  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R�*!��������؉�����u!hpj h�  h�j�3������u̃����� uI��0���    j h�  h�h�hp�*����ǅ����������T����<1���������  �'  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��D�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Yh�  h�j��d���]  P����������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�E���E�M�Q��A��������������  ������ |������d}ǅH���   �
ǅH���    ��H��������������� u!h 	j h  h�j�������u̃����� uI�/���    j h  h�h�h 	�c(����ǅ����������T����/����������  ��@���t!h0j h  h�j�������u̋����������������������������������������Q��A���������������T����#��P��h���Q��d���R��D���P��P���Q������R������P��AQ�ܑ�Ѓ���������   t.��d��� u%��T�������P������P��AQ�ܑ�Ѓ���D�����gu2������%�   u%��T������P������Q��AR�ܑ�Ѓ����������-u!��������   ��������������������������Q�@�����������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ������%�   t&�0   f��������4�����Qf������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  �%  ������ u�EP�������������������  ������ |������d}ǅD���   �
ǅD���    ��D��������������� u!h 	j h�  h�j�{������u̃����� uI�	,���    j h�  h�h�h 	�S%����ǅ����������T����,����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�`��������؉�����u!h�j h�  h�j�i������u̃����� uI��*���    j h�  h�h�h��A$����ǅ����������T����r+����������  �]  �1��������������������������Q������������������  ��������   �%  ������ u�EP��������������������  ������ |������d}ǅ@���   �
ǅ@���    ��@��������������� u!h 	j h�  h�j�D������u̃����� uI��)���    j h�  h�h�h 	�#����ǅ����������T����M*���������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�)��������؉�|���u!h�j h�  h�j�2������u̃�|��� uI��(���    j h�  h�h�h��
"����ǅ����������T����;)���������  �&  �1����������������x�����x���Q��������������������  �������� �e  ��������@�)  ������ u�MQ��%��������������������  ������ |������d}ǅ<���   �
ǅ<���    ��<�����t�����t��� u!h 	j h�  h�j��������u̃�t��� uI�'���    j h�  h�h�h 	�� ����ǅ����������T����(���������_  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q����������؉�p���u!h�j h�  h�j��������u̃�p��� uI�{&���    j h�  h�h�h�������ǅ����������T�����&���������M  ��  �3����������������l�����l���R��#�������������������(  ������ u!�EP�#���������������������  ������ |������d}ǅ8���   �
ǅ8���    ��8�����h�����h��� u!h 	j h�  h�j��������u̃�h��� uI�b%���    j h�  h�h�h 	�����ǅ����������T�����%���������4  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P���������؉�d���u!h�j h�  h�j��
������u̃�d��� uI�P$���    j h�  h�h�h������ǅ����������T�����$���������"  �  �5����������������`�����`���Q�!��������������������Z  ��������@�'  ������ u�EP�f!�������������������  ������ |������d}ǅ4���   �
ǅ4���    ��4�����\�����\��� u!h 	j h  h�j�	������u̃�\��� uI�)#���    j h  h�h�h 	�s����ǅ����������T����#����������
  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P���������؉�X���u!h�j h  h�j�������u̃�X��� uI�"���    j h  h�h�h��a����ǅ����������T����"����������	  �}  �2����������������T�����T���Q�f������������������$  ������ u�UR�?����3ɉ�������������  ������ |������d}ǅ0���   �
ǅ0���    ��0�����P�����P��� u!h 	j h0  h�j�s������u̃�P��� uI�!���    j h0  h�h�h 	�K����ǅ����������T����|!����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�X��������؉�L���u!h�j h4  h�j�a������u̃�L��� uI�����    j h4  h�h�h��9����ǅ����������T����j ����������  �U  �3����������������H�����H���R�>����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ��������������d��� }ǅd���   �%�����������������d���   ~
ǅd���   �����������u
ǅ����    ��O�����������d�����d�������d������������������   �������RP������P������Q�m����0�������������RP������R������P����������������������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�k  ��l��� �:  ��������@tj��������   t�-   f������ǅ����   �D��������t�+   f������ǅ����   �!��������t�    f������ǅ����   ������+�����+�������D�����������u��L���Q�UR��D���Pj ��  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��D���Qj0�  �������� ��   ������ ��   ��������@�����������<�����<�����<�������<�������   ��T������P��T����y��� ���   Q��@���R��<���P�������8�����8��� ǅL��������2��L���Q�UR��<���P�E  ����@����8�����@����`����(��|���R��L���P�MQ������R������P��  ����L��� |'��������t��L���R�EP��D���Qj �T  �������� tj������R�����ǅ����    ������8��� t��8���tǅ,���    �
ǅ,���   ��,�����4�����4��� u!hhj h�  h�j�� ������u̃�4��� uI�^���    j h�  h�h�hh�����ǅ����������T��������������0  �������  ��@��� ��  ǅ����    ���������������������;�x�����  ����������������(�����(�������(�����(�����   ��(����$���
���������E�������MQ�4�����_  ���������E�������MQ������;  ���������E�������MQ������  ���������E�������MQ�������   ���������E�������MQ�������   ���������E�������MQ�g�����������������   3�tǅ$���   �
ǅ$���    ��$�����0�����0��� u!h�j h.	  h�j���������u̃�0��� uF�R���    j h.	  h�h�h������ǅ����������T��������������'�����#�����L�����������T�������������M�3��A�����]Ë��{
�{
&|
�|
�
�
d�
փ
�|
�|
p|
_|
�|
�|
 �I ݂
��
��
��
у
 ��
�
��
g�
�
7�
0�
0�
�
��
]�
��
N�
s�
A�
   	
��
"�
F�
j�
��
�
��
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U��j�h6h�d�    P���SVW��A1E�3�P�E�d�    3��} ���E܃}� uhlj j3h�j�t�������u̃}� u-����    j j3h�h�hl�R �������  �M�U�U�E�P�Y������E�    �M�Q�UR� ����f�E��E������   ��E�P��������f�E��M�d�    Y_^[��]����������������������������������������������������������������������������̋�U���8��A3ŉE�V�E�H��@�d  �UR�q��������t@�EP�`��������t/�MQ�O����������UR�>�������������E���E�B�E�H$�����у�tj�EP���������t@�MQ����������t/�UR������������EP���������������E���E�B�M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ�������  �(  �UR�5��������t@�EP�$��������t/�MQ�����������UR��������������E���E�B�E��H��   ��   �URj�E�P�M�Q�������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R�������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP�.�����^�M�3�������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�p�����]��������̋�U���8�EP�M�����3Ƀ} ���M�}� uh0�j j4h�j��������u̃}� u=����    j j4h�h�h0��`������E�����M�����E��  3��} ���E��}� uh��j j5h�j��������u̃}� u=����    j j5h�h�h����������E�����M��$���E��   �M�� �����z u"�EP�MQ�������EԍM������E��x�b�U��E̍M������P�M�Q��������E��U���U�E��MȍM�����P�U�R�������E��E���E�}� t�M�;M�t��U�+U��UЍM��w���EЋ�]����������������������������������������������������������������������������������������������������������̋�U����E��M��U��E���E��A|�}�Z	�M��� �M��U��E��M��U���U��A|�}�Z	�E��� �E��}� t�M�;M�t��E�+E���]������������������������������̋�U����=�m ��   3��} ���E��}� uh0�j jbh�j���������u̃}� u0�r����    j jbh�h(h0������������   3҃} �U��}� uh��j jch�j�{�������u̃}� u-�����    j jch�h(h���Y����������&�MQ�UR��������j �EP�MQ���������]������������������������������������������������������������������������̋�U���@�} �!  �EP�M�����3Ƀ} ���M�}� uh0�j j;h�j��������u̃}� u=�����    j j;h�hhh0��f������E�����M������E��  3��} ���E��}� uh��j j<h�j��������u̃}� u=�����    j j<h�hhh����������E�����M��*����E��1  ����;U����E�uh@j j=h�j��������u̃}� u=�3����    j j=h�hhh@�������E�����M������E��   �M�������z u)�EP�MQ�UR��������E̍M������E��   �m�E��MčM��q���P�U�R�Z������E��E���E�M��U��M��G���P�E�P�0������E��M���M�U���Ut�}� t�E�;E�t��M�+M��MȍM�������E��3���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����=�m �Y  3��} ���E��}� u!h0�j h�   h�j��������u̃}� u3�O����    j h�   h�h h0������������  3҃} �U��}� u!h��j h�   h�j�R�������u̃}� u3������    j h�   h�h h���-����������   ����;M҃��U�u!h@j h�   h�j���������u̃}� u0�w����    j h�   h�h h@������������.�MQ�UR�EP�[�������j �MQ�UR�EP���������]��������������������������������������������������������������������������������������������������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   ��}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q���_^��]� ���������������������̋�U��Q�M��E�� D�M��A    �U��B �E���]����������������������̋�U��Q�M��M��B����E��t�M�Q�c������E���]� �����������������̋�U��Q�M��E�� D�M��A    �U��B �E�Q�M��Z����E���]� ���������������������̋�U��Q�M��E�� D�M��U��A�M��A �E���]� ������������������̋�U��Q�M��E�� D�M��A    �U��B �EP�M��:����E���]� �����������������������̋�U��Q�M��E�;Et0�M��"����M�Q��t�E�HQ�M��x�����U��E�H�J�E���]� ���������������������̋�U��Q�M��E�� D�M��������]������������������̋�U����M��E��x t�M��Q�U���E�P�E���]�������������������̋�U����M��} tK�EP�8��������E��M�Q�+������U��B�E��x t�MQ�U�R�E��HQ�f������U��B��]� �����������������������������̋�U��Q�M��E��H��t�U��BP�������M��A    �U��B ��]������������������������̋�U��Q�M��EP�M������M��l�E���]� ��������̋�U��Q�M��M��%����E��t�M�Q�s������E���]� �����������������̋�U��Q�M��EP�M������M��l�E���]� ��������̋�U��Q�M��E�� l�M��������]������������������̋�U��Q�M��EP�M������M��|�E���]� ��������̋�U��Q�M��M�������E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M�������M��|�E���]� ��������̋�U��Q�M��E�� |�M��	�����]������������������̋�U��Q�M��EP�M������M����E���]� ��������̋�U��Q�M��M������E��t�M�Q��������E���]� �����������������̋�U��Q�M��EP�M������M����E���]� ��������̋�U��Q�M��E�� ��M�������]������������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���������������������������̋�U��j j jj jh   @h�����V]����������̋�U��=�V�t�=�V�t��VP��]�����������̋�U��j�h86h�d�    P���SVW��A1E�3�P�E�d�    �E�����3��} ���E��}� uh��j j.h�j��������u̃}� u+�����    j j.h�h�h���k���������W�U�B��@t�M�A    �=�UR�c������E�    �EP�w������E��E������   ��MQ�������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U����E�����3��} ���E�}� uhlj jYh�j�g�������u̃}� u.������    j jYh�h4hl�E���������   �U�U��E��H��   ta�U�R�i������E��E�P�������M�Q������P���������}	�E������$�U��z tj�E��HQ�5������U��B    �E��@    �E���]�����������������������������������������������������������������������̋�U��j�hX6h�d�    P���SVW��A1E�3�P�E�d�    �}�u������ 	   ����  �} |�E;<�s	�E�   ��E�    �M؉M��}� uh(j j,h�j���������u̃}� u.�a���� 	   j j,h�h�h(����������;  �E���M���������D
������؉E�uhXj j-h�j�U�������u̃}� u.������ 	   j j-h�h�hX�3����������   �UR�h������E�    �E���M���������D
��t;�MQ�������P����u�$��E���E�    �}� u�>������U��J���� 	   �E�����3�uhX�j jEh�j��������u��E������   ��UR�������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�   ��]�������������������̋�U���$�} t�E�M�3҃} �U�}� uhLj j^h�j�P�������u̃}� u-������    j j^h�h�hL�.�����3��'  �} t�}|�}$~	�E�    ��E�   �M��M�}� uh`j j_h�j���������u̃}� u-�b����    j j_h�h�h`������3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q���������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R�V�������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q��������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q��������E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4������ "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�X�����]�������������������̋�U��j�EP�MQ�UR�(�����]�������������������̋�U��j�EP�MQ�UR�������]�������������������̋�U��� �} uh`�j jdh�j�J�������u̋M�M��U�R�A������E��E��H��   u&����� 	   �U��B�� �M��A���  �c  �/�U��B��@t$����� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6������ 9E�t������@9E�u�M�Q���������u�U�R�E������E��H��  �  �U��E��
+Hy!hP�j h�   h�j���������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�������E��s�}��t!�}��t�M����U���������U���E�B�E��H�� t9jj j �U�R��������E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q�P������E�U�;U�t�E��H�� �U��J���  ��E%��  ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̋�U��j�hx6h�d�    P���SVW��A1E�3�P�E�d�    �}�u�7����     ����� 	   ����  �} |�E;<�s	�E�   ��E�    �M؉M��}� uh��j j.hPj���������u̃}� u9������     �K���� 	   j j.hPh<h������������  �E���M���������D
������؉E�uh�j j/hPj�?�������u̃}� u9�B����     ������ 	   j j/hPh<h�����������   �UR�G������E�    �E���M���������D
��t�MQ��������E��4�S���� 	   �E�����3�uhX�j j9hPj��������u��E������   ��MQ�������ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QV�EP���������t]�}u������   ��u�}u(����HD��tj�q�������j�e�����;�t�UR�U�����P����t	�E�    �	�$��E��EP�0������M���U���������D �}� t�M�Q����������3�^��]����������������������������������������������������̋�U��} uh8j j.h�j��������u̋M�Q��   tK�E�H��t@j�U�BP��������M�Q�������E�P�M�    �U�B    �E�@    ]��������������������������������������������̋�U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%ؑ�%ܑ�%���%��%��%��%��%���%���%���% ��%��%��%��%��%��%��%��% ��%$��%(��%,��%0��%4��%8��%<��%@��%D��%H��%L��%P��%T��%X��%\��%`��%d��%h��%l��%p��%t��%x��%|��%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%Ē�%Ȓ�%̒�%В�%Ԓ�%ؒ�%ܒ�%���%��%��%��%��%���%���%���% ��%��%��%��%��%��%����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍M������T$�B�J�3�誴���(/����������������̡Dm����DmËT$�B�J�3��t�����/�Y�������������������������̍M������T$�B�J�3��:�����0����������������̋T$�B�J�3������l4�������������������������̍M��>����T$�B�J�3��ڳ����4����������������̍M������T$�B�J�3�誳����4�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������PX�i���h@薩����_^[���   ;�������]������������������������U����   SVW��@����0   ������j �]貭��_^[���   ;��ĸ����]������������������̋�U��Q3��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������PX�L���_^[���   ;��V�����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         p�
��
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �8��լ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            -�:�                                                                                                                                                                                                                                                                    ߶                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �u=P       {   � �r          �p@              @             �o@                    PointCount:               �?        c:\program files\maxon\cinema 4d r13\plugins\drawtext tag_r13\source\drawtext tag.cpp                   PolyCount:      tsimpletag      myicon.png       Ҡ@�"���ʼG�m������C����H�c����~�����                    P#� �"���ʼ�m������C����H�y���������                    h$� �"���ʼ�m������C����H�y����                IDM_NEU     SDK Test    IDS_EDITOR_PLUGINS      PLUGIN_CMD_1000472      M_EDITOR    C4DSDK - Edit Image Hook:       -plugincrash    -SDK executed:-)       -SDK    -SDK is here :-)       -help   --help  res c:\program files\maxon\cinema 4d r13\resource\_api\c4d_memory.cpp               c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp                  %s      c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h                c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp                 #   ���        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp             �ǰ    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp                 ���    � ��    � ��    � ��    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_string.cpp               no baselist      B   KB  MB           �@     GB c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp                c:\program files\maxon\cinema 4d r13\resource\_api\ge_sort.cpp              U�T!��        f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c                            f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c             Unknown Runtime Check Error
       Stack memory around _alloca was corrupted
         A local variable was used before it was initialized
           Stack memory was corrupted
        A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                �E0DD�C�CtC                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                  Run-Time Check Failure #%d - %s         Unknown Module Name     Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s                   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                           Stack corrupted near unknown variable               Stack area around _alloca memory reserved by this function is corrupted
                %s%s%s%s    >   
   %s%s%p%s%ld%s%d%s           Stack area around _alloca memory reserved by this function is corrupted                 
Address: 0x    
Size:      
Allocation number within this function:            
Data: <    wsprintfA   u s e r 3 2 . d l l         %.2X    A variable is being used without being initialized.             Stack around _alloca corrupted          Local variable used before initialization           Stack memory corruption     Cast to smaller type causing loss of data           Stack pointer corruption        K�J�J�J\J    f:\dd\vctools\crt_bld\self_x86\crt\prebuild\misc\i386\chkesp.c                  The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                       _ s e t d e f a u l t p r e c i s i o n                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c                         s i z e I n B y t e s   >   0           _ c f t o e _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c                         b u f   ! =   N U L L       e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                           _ c f t o e 2 _ l           s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o a _ l         _ c f t o f _ l         _ c f t o f 2 _ l       _ c f t o g _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p                             p N o d e - > _ N e x t   ! =   N U L L                 s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                 f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c           FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    K E R N E L 3 2 . D L L         Client  Ignore  CRT Normal  Free    (T TTTT    Error: memory allocation: bad memory block type.
           Invalid allocation size: %Iu bytes.
        Client hook allocation failure.
        Client hook allocation failure at file %hs line %d.
            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c                         _ C r t C h e c k M e m o r y ( )           _ p F i r s t B l o c k   = =   p O l d B l o c k               _ p L a s t B l o c k   = =   p O l d B l o c k             f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       Error: possible heap corruption at or near 0x%p                 p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Client hook re-allocation failure.
         Client hook re-allocation failure at file %hs line %d.
             _ e x p a n d _ d b g       p U s e r D a t a   ! =   N U L L           _ p F i r s t B l o c k   = =   p H e a d           _ p L a s t B l o c k   = =   p H e a d             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                                 HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()                _ m s i z e _ d b g         %hs located at 0x%p is %Iu bytes long.
             %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
                   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 DAMAGED     _heapchk fails with unknown return value!
          _heapchk fails with _HEAPBADPTR.
       _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADBEGIN.
         _ C r t S e t D b g F l a g             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t D o F o r A l l C l i e n t O b j e c t s               p f n   ! =   N U L L       Bad memory block found at 0x%p.
        Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              _ C r t M e m C h e c k p o i n t           s t a t e   ! =   N U L L           n e w S t a t e   ! =   N U L L         o l d S t a t e   ! =   N U L L         _ C r t M e m D i f f e r e n c e           Object dump complete.
      crt block at 0x%p, subtype %x, %Iu bytes long.
             normal block at 0x%p, %Iu bytes long.
          client block at 0x%p, subtype %x, %Iu bytes long.
              {%ld}   %hs(%d) :       #File Error#(%d) :      Dumping objects ->
      Data: <%s> %s
     ( * _ e r r n o ( ) )       _ p r i n t M e m B l o c k D a t a             Detected memory leaks!
     Total allocations: %Id bytes.
          Largest number used: %Id bytes.
        %Id bytes in %Id %hs Blocks.
       _ C r t M e m D u m p S t a t i s t i c s           o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g               Damage before 0x%p which was allocated by aligned routine
                  The block at 0x%p was not allocated by _aligned routines, use realloc()                 The block at 0x%p was not allocated by _aligned routines, use free()                _ a l i g n e d _ m s i z e _ d b g             m e m b l o c k   ! =   N U L L         CorExitProcess      m s c o r e e . d l l       _ w p g m p t r   ! =   N U L L         _ g e t _ w p g m p t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 d a t . c                         p V a l u e   ! =   N U L L         _ p g m p t r   ! =   N U L L           _ g e t _ p g m p t r       f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c             s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               _ s e t e n v p             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c            f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c            f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c          f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h e a p i n i t . c                       _ c r t h e a p           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                                      H_�_        ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                 _ v s n p r i n t f _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c                       ( f o r m a t   ! =   N U L L )         r u n t i m e   e r r o r            
     T L O S S   e r r o r  
           S I N G   e r r o r  
         D O M A I N   e r r o r  
             R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                            �x   �x	   x
   �w   Hw   �v   �v    v   �u   @u   �t   @t   �s   �s   �r    (r!   �ox   �oy   �oz   lo�   do�   @o                                        M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             
 
     w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                               . . .       w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           < p r o g r a m   n a m e   u n k n o w n >             w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                             R u n t i m e   E r r o r ! 
 
 P r o g r a m :                     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     _ N M S G _ W R I T E           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c                         s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         _ _ g e t l o c a l e i n f o               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t h e l p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\inithelp.c           M S P D B 1 0 0 . D L L     M S V C R 1 0 0 D . d l l               r   PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y                 S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S                       RegCloseKey     RegQueryValueExW    RegOpenKeyExW   A D V A P I 3 2 . D L L         D L L       M S P D B 1 0 0         ... Assertion Failed    Error   Warning     ��؁ā    f:\dd\vctools\crt_bld\self_x86\crt\src\dbgrpt.c             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       p f n N e w H o o k   ! =   N U L L             _ C r t S e t R e p o r t H o o k 2                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c                           m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           Microsoft Visual C++ Debug Library          _CrtDbgReport: String too long or IO Error          s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                     Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)                    
Module:    
File:      
Line:      

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.                              m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                 <program name unknown>      s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         _ _ c r t M e s s a g e W i n d o w A           A s s e r t i o n   F a i l e d         E r r o r       W a r n i n g       d�T�,�    _ C r t S e t R e p o r t H o o k W 2           M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y                     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )                                     
 M o d u l e :         
 F i l e :         
 L i n e :         E x p r e s s i o n :               
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                     w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       _ _ c r t M e s s a g e W i n d o w W           _ c o n t r o l f p _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c                           ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c                       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )                                                                                         H H : m m : s s         d d d d ,   M M M M   d d ,   y y y y           M M / d d / y y         P M     A M     D e c e m b e r         N o v e m b e r         O c t o b e r       S e p t e m b e r       A u g u s t     J u l y     J u n e     A p r i l       M a r c h       F e b r u a r y         J a n u a r y       D e c       N o v       O c t       S e p       A u g       J u l       J u n       M a y       A p r       M a r       F e b       J a n       S a t u r d a y         F r i d a y     T h u r s d a y         W e d n e s d a y       T u e s d a y       M o n d a y     S u n d a y     S a t       F r i       T h u       W e d       T u e       M o n       S u n       HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun p f l t   ! =   N U L L             s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           _ f p t o s t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c                       _ g e t _ e r r n o             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d o s m a p . c                       _ g e t _ d o s e r r n o           s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                     _ f l t o u t 2             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c                         _ s e t _ o u t p u t _ f o r m a t             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t f o r m a t . c                               ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                   ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               B u f f e r   i s   t o o   s m a l l           ( ( ( _ S r c ) ) )   ! =   N U L L             s t r c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                     f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c           Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete      new    __unaligned     __restrict      __ptr64     __eabi  __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(    ������ؠ̠Ġ�������K������|�x�t�p�l�h�\�X�T�P�L�H�D�@�<�8�4�0�,�(�$� �������� �������������ԟȟ��������p�L�(��������p�H� ��Н��������p�h�\�H�(��Ԝ��x�D�$���Л��h�D��K,���̚��                                                                                CV:     ::  '   `   generic-type-   template-parameter-     ''  `anonymous namespace'       `non-type-template-parameter        `template-parameter     void    NULL    extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{        }'  }'  )   void    std::nullptr_t      volatile    ,<ellipsis>     ,...    <ellipsis>       throw(      volatile   const   signed      unsigned    UNKNOWN     __w64   wchar_t     <unknown>   __int128    __int64     __int32     __int16     __int8  bool    double  long    float   long    int short   char    enum    cointerface     coclass     class   struct      union   `unknown ecsu'      int     short   char    const   volatile    cli::pin_ptr<   cli::array<     )[  {flat}  s   {for    ������    ����@�    ��;���    ������    ��}�ө     ??     �|���    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h a n d l e r . c p p                         p n h   = =   0         _ e x p a n d _ b a s e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c                       p B l o c k   ! =   N U L L         ( s t r i n g   ! =   N U L L )         s p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c                         ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6             s i g n a l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c                       ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f:\dd\vctools\crt_bld\self_x86\crt\src\winsig.c             r a i s e       SystemFunction036           ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       r a n d _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r a n d _ s . c                       _ R a n d o m V a l u e   ! =   N U L L             ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c                         s t r   ! =   N U L L       ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c             ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 ( c h   ! =   _ T ( ' \ 0 ' ) )         (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       _ o u t p u t _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c                       ( s t r e a m   ! =   N U L L )         _ s e t _ e r r o r _ m o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c                         ( " I n v a l i d   e r r o r _ m o d e " ,   0 )               GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L             ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               w c s c a t _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                     w c s n c p y _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l                         w c s c p y _ s         s t r n c p y _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h                           ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                   _ w m a k e p a t h _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t m a k e p a t h _ s . i n l                         ( L " I n v a l i d   p a r a m e t e r " ,   0 )               _ w s p l i t p a t h _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t s p l i t p a t h _ s . i n l                           ( ( ( _ P a t h ) ) )   ! =   N U L L           f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t M o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c                         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   _ C r t S e t R e p o r t F i l e               _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       %s(%d) : %s         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed!       Assertion failed:           s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   , Line      <file unknown>      Second Chance Assertion Failed: File            _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t A           w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               _CrtDbgReport: String too long or Invalid characters in String                  s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       % s ( % d )   :   % s       w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                 w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d !           A s s e r t i o n   f a i l e d :                   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 
   ,   L i n e         < f i l e   u n k n o w n >             S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t W           GetUserObjectInformationA       MessageBoxA     s i z e I n B y t e s   > =   c o u n t             s r c   ! =   N U L L       m e m c p y _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c                       d s t   ! =   N U L L       _ s w p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s w p r i n t f . c                            _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                         _ s e t _ c o n t r o l f p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                             LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL  p�    c�`��H�T��H��D��Hz�4��H��(��H��                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         _ c o n f i g t h r e a d l o c a l e           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t l o c a l . c                       ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                       f:\dd\vctools\crt_bld\self_x86\crt\src\setlocal.c           s e t l o c a l e       L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     s t r n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ s e t l o c a l e _ n o l o c k           ;   =;  s t r c p y _ s ( p c h   +   s i z e o f ( i n t ) ,   c c h   -   s i z e o f ( i n t ) ,   l c t e m p )                         _ s e t l o c a l e _ s e t _ c a t             s t r c a t _ s ( p c h ,   c c h ,   " ; " )               _ s e t l o c a l e _ g e t _ a l l             s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   s t r n c p y _ s ( c a c h e i n ,   c a c h e i n S i z e ,   s o u r c e ,   c h a r a c t e r s I n S o u r c e   +   1 )                               C   s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   " C " )                 _ e x p a n d l o c a l e           s t r c a t _ s ( o u t s t r ,   s i z e I n B y t e s ,   (   * ( c h a r   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                           _ s t r c a t s             s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                               s t r n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   l o c a l e ,   l e n )                                             s t r n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                           _., s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & l o c a l e [ 1 ] ,   1 6 - 1 )                                             _ _ l c _ s t r t o l c         .   _   s t r c p y _ s ( l o c a l e ,   s i z e I n B y t e s ,   ( c h a r   * ) n a m e s - > s z L a n g u a g e )                         _ _ l c _ l c t o s t r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t t i m e . c                       p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                   f:\dd\vctools\crt_bld\self_x86\crt\src\inittime.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t n u m . c                         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initnum.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t m o n . c                         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initmon.c                                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                            _ _ s t r g t o l d 1 2 _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l                             _ L o c a l e   ! =   N U L L           1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 $ I 1 0 _ O U T P U T       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c                             _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r           _ v s n p r i n t f _ h e l p e r           ( " B u f f e r   t o o   s m a l l " ,   0 )               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   _ v s p r i n t f _ s _ l           f o r m a t   ! =   N U L L         _ v s n p r i n t f _ s _ l         ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   ( _ o s f i l e ( f h )   &   F O P E N )           _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c                       ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c                     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )               ( ( c n t   &   1 )   = =   0 )         _ w r i t e _ n o l o c k           ( b u f   ! =   N U L L )           f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c                         _ i s a t t y           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c          _ f i l e n o       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c                       p r i n t f         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p r i n t f . c                       _ w c t o m b _ s _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c                       s i z e I n B y t e s   < =   I N T _ M A X             _ m b s t o w c s _ l _ h e l p e r                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c                       s   ! =   N U L L       r e t s i z e   < =   s i z e I n W o r d s             b u f f e r S i z e   < =   I N T _ M A X           _ m b s t o w c s _ s _ l           ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                               s t r c a t _ s         l e n g t h   <   s i z e I n T C h a r s           2   < =   r a d i x   & &   r a d i x   < =   3 6               s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   s i z e I n T C h a r s   >   0         x t o a _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c                       x 6 4 t o a _ s         _ w c s t o m b s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c                       p w c s   ! =   N U L L         s i z e I n B y t e s   >   r e t s i z e           _ w c s t o m b s _ s _ l           ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               _ v s w p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c                       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s w p r i n t f _ s _ l         _ v s n w p r i n t f _ s _ l           x t o w _ s     x 6 4 t o w _ s         _ w o u t p u t _ l         _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             p l o c i - > c t y p e 1 _ r e f c o u n t   >   0                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t c t y p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\initctyp.c           united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american    ��ENU ��ENU ��ENU ��ENA ��NLB ��ENC ��ZHH |�ZHI p�CHS \�ZHH D�CHS ,�ZHI �CHT �NLB ��ENU ��ENA ��ENL ��ENC ��ENB ��ENI ��ENJ p�ENZ T�ENS 4�ENT $�ENG �ENU �ENU ��FRB ��FRC ��FRL ��FRS ��DEA ��DEC p�DEL `�DES P�ENI @�ITS 4�NOR  �NOR �NON ��PTB ��ESS ��ESB ��ESL ��ESO ��ESC d�ESD P�ESF 8�ESE  �ESG �ESH ��ESM ��ESN ��ESI ��ESA ��ESZ ��ESR |�ESU h�ESY P�ESV <�SVF 4�DES 0�ENG ,�ENU (�ENU                                                                                                         �USA �GBR �CHN  �CZE ��GBR ��GBR ��NLD ��HKG ��NZL ��NZL ��CHN ��CHN ��PRI ��SVK x�ZAF h�KOR X�ZAF H�KOR 0�TTO 0�GBR �GBR �USA ,�USA                                     6-    Norwegian-Nynorsk           s t r c p y _ s ( l p O u t S t r - > s z L a n g u a g e ,   ( s i z e o f ( l p O u t S t r - > s z L a n g u a g e )   /   s i z e o f ( l p O u t S t r - > s z L a n g u a g e [ 0 ] ) ) ,   " N o r w e g i a n - N y n o r s k " )                                                   _ _ g e t _ q u a l i f i e d _ l o c a l e                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t q l o c . c                         OCP ACP ܾbad exception   �!R���        i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                   s t r t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o l . c                       n p t r   ! =   N U L L         s t r t o x q       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o q . c                           ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 _ o u t p u t _ p _ l           ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f:\dd\vctools\crt_bld\self_x86\crt\src\osfinfo.c            _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c                           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                             f:\dd\vctools\crt_bld\self_x86\crt\src\_sftbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ s f t b u f . c                         f l a g   = =   0   | |   f l a g   = =   1             v p r i n t f _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v p r i n t f . c                         _ w o u t p u t _ s _ l         _ w o u t p u t _ p _ l         f p u t w c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t w c . c                       ( s t r   ! =   N U L L )           _ s t r i c m p _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r i c m p . c                         _ s t r i c m p         c o u n t   < =   I N T _ M A X         _ s t r n i c m p _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c m p . c                       _ s t r n i c m p       csm�               �                H"����    Unknown exception       `"����    �"ҥ��    #s���    C O N O U T $       f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c                       _ f c l o s e _ n o l o c k         ( _ o s f i l e ( f i l e d e s )   &   F O P E N )             _ c o m m i t           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c                           ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         w c s t o x l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o l . c                       _ c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c                     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c                       s t r e a m   ! =   N U L L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         RSDS���v3/�K��V��)   C:\Program Files\MAXON\CINEMA 4D R13\plugins\DrawText Tag_R13\obj\DrawText Tag_R13_Win32_Debug.pdb                                                                                                                                                                                                                                                                                                      @8               L    `��    @       ����    @   8         @       ����    @   �                   �    ��    <@       ����    @   �                       �    X@        ����    @   4                   H                     @�                <@�                X@4                �@�               �    �    �@        ����    @   �                    �@                     ( L     �@       ����    @            �@        ����    @   p                    �     L                 �@p                 A�                �     �     A        ����    @   �                     0A!               (!    0!    0A        ����    @   !                    pAl!               �!    �!    pA        ����    @   l!                    �R�!               �!    �!"    �R       ����    @   �!        �R        ����    @   ,"                   @"    "                �R,"                hVx"               �"    �""    hV       ����    @   x"                    �V�"               �"    �""    �V       ����    @   �"                    �V0#               D#    T#�""    �V       ����    @   0#                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ����    ����    ����    W�    ����    ����    ����e���    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����v�|�    ����    ����    ����    �%    ����    ����    ����    �'    ����    ����    ����    >)    ����    ����    ����    �+    ����    ����    ����    �,    ����    ����    ����    �1����    	2        ����    ����    ����    �4����    e5        ����    ����    ����    <    ����    ����    ����    R?    ����    ����    ����    I    ����    ����    ����    J    ����    ����    ����    FR    ����    ����    ����    �S    ����    ����    ����    �X    ����    ����    ����    V[    ����    ����    ����    �\    ����    ����    ����    _    ����    ����    ����    b    ����    ����    ����    jh    ����    ����    ����    �}    ����    ����    ����    ��    ����    ����    ����    &�    ����    ����    ����    Q�    ����    ����    ����    �    ����0�
"�    /                           ����    ����    ����    ��    ����    ����    ����    �	    ����    x���    ����    �    ����    x���    ����    c    ����`�
"�   �/                           ����    ����    ��������    ����    ����    ��������    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    Y�    ����    ����    ����    :�    ������
"�   �0                           ����    ����    ����    �>        �=        ����    |��    ����    7J        �G        ����    ����    ����    �e    ����    ����    ����    �f����    g        ����    ����    ����    bk����    �k        ����    ����    ����    Gn        Lm        n            ����    ����    ����    T�    ����    ����    ����    ? 	    ����    ����    ����    �	    ����    ����    ����gt	�t	        ��    �2       �2�2        �R    ����       �        �R    ����       �        ����    ����    ����    }�	    M�	Z�	        ����    ����    ����    ��	    ��	�	        ����    ����    ����&�	,�	    ����    ����    ����շ	۷	    ����    ����    ����ø	θ	    ����    ����    ����{�	��	    ����    ����    �����	,�	    ����    ����    ������	��	    ����    ����    ����h�	u�	    @           ��	����    ����                  84"�   H4   X4                       ���� �
"�   �4                           ����0�
"�   �4                           ����    ����    ����    �B
        sA
        ����    ����    ����    3I
    ����    ����    ����    �J
    ����    ����    ����    "L
    ����    ����    ����    �P
    ����    ����    ����    �Q
    ����    ����    ����    �T
        �T
        ����    ����    ����    �X
    ����    ����    ����    �
    ����    ����    ����    ��
    ����    ����    ����    ��
    ����    ����    ����    |�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �u=P    "9          9 9  9 ˬ 79   DrawText Tag_R13.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 V   �B    .?AVSimpleTag@@     �B    .?AVTagData@@       �B    .?AVNodeData@@      �B    .?AVBaseData@@      �   �   �   �   �  �  B  8   ^  �  �B    .?AVGeToolDynArray@@        -   �B    .?AVGeToolDynArraySort@@        �B    .?AVGeSortAndSearch@@       �B    .?AVGeToolList2D@@      �B    .?AVGeToolNode2D@@         Q   �   u�  s�              �B    .?AVtype_info@@         N�@���D                           1�1�1�1�1�1�1�1�1�1�        ��������       ����   ��������        �����
                                                                         ���{                                                                                                                                                                                                                                                                                                                                    abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     hB�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ����C   ������������������|�p�d�\�P�L�H�D�@�<�8�4�0�,�(�$� ��� ���<�����ԓȓ������������x�	         l�`�T�H�<�0�$����ؒ����������t�h�\�P�D�8�,� �����ܑ̑��\�������|�h�P�8�0�(����Ȑ                                                                                                                                                                   �H            �H            �H            �H            �H                              �N        0���8��H                                            HJHJhB                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��            ��|�    ����         ������������        4�    .   .   �N�m�m�m�m�m�m�m�m�m�N�m�m�m�m�m�m�m�N                    0�2�       ���5      @   �  �   ����                          �                     q     q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �D        � 0                .              �B    .?AVbad_exception@std@@         �B    .?AVexception@std@@                      �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                            �B    .?AVbad_cast@std@@      �B    .?AVbad_typeid@std@@        �B    .?AV__non_rtti_object@std@@                 ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (�         d� ؑ                     �� �� �� �� Г � �� � "� .� @� P� l� x� �� �� �� �� ʔ ڔ � � � &� 6� D� V� f� �� �� �� ƕ ܕ �� � � ,� F� V� l� �� �� �� ʖ � �� 
� � (� 4� F� V� d� n� z� �� �� �� ȗ ؗ � � �� � .� D� Z� j� �� �� �� �� Ę ֘ � �� � $� 4� B� P�                                                                                                             �� �� �� �� Г � �� � "� .� @� P� l� x� �� �� �� �� ʔ ڔ � � � &� 6� D� V� f� �� �� �� ƕ ܕ �� � � ,� F� V� l� �� �� �� ʖ � �� 
� � (� 4� F� V� d� n� z� �� �� �� ȗ ؗ � � �� � .� D� Z� j� �� �� �� �� Ę ֘ � �� � $� 4� B� P�                                                                                                             �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer WideCharToMultiByte  IsDebuggerPresent gMultiByteToWideChar �RaiseException  MlstrlenA  EGetProcAddress  ?LoadLibraryW  IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  GetLastError  �InterlockedDecrement  �GetCurrentThread  �HeapValidate  �IsBadReadPtr  ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter GetModuleFileNameW  %WriteFile GetLocaleInfoW  �HeapFree  �HeapAlloc JGetProcessHeap  �VirtualQuery  bFreeLibrary hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage � EnterCriticalSection  9LeaveCriticalSection   FatalAppExitA RtlUnwind �HeapReAlloc �HeapSize  �HeapQueryInformation  -SetConsoleCtrlHandler �InterlockedExchange �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -LCMapStringW  iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  GetLocaleInfoA  IsValidLocale EnumSystemLocalesA  �GetUserDefaultLCID  �SetStdHandle  � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �    �:];v;�;<�<=�>�?�? � H   0#0\0a0j0�0�0�0�0�0&1+141R1�:�;�;�;<<<A<L<j<�<�<�<�<
===8=     (   7,787D7P7\7h7t7�7�7�7�7�7�7�?�?  D   [0�01�1g2;3�374j4�4�45�56�67�7/89�9$;=�=�=>W>|>�>�?�?   L   P0 1�2�4�4Q5�5�5�596�6Y7|7�7�8r9�9�:�:�: ;
;�;Q<o<�<�<�<=w=�>??   0 T   m3w3�3�3�3�3�3�3�3�3�3�3�3�3�344545@5,6R9W9�9&:�:
;z;�;�<�<�=>A>�>?�?�? @ X   \0�0�0%1�12p2�203o3�3m4�4�4�4Z5�5�56]6b6�6f7�7F8�89�9::�:h;�;�<==>�>?�? P <   0�01�12�23�3C4�4+5�526�6+7�788�8�9
:�:;;�;�;�; ` ,   L0Q0k0p0H1M1?4�4G5�5;6�6�;�;<<�<   p T   �1�1�1�2�2/3�3�3�3�3x4}4�4?5d5p5|5�5h6�6o7�7_8�899:�:g;�;_<�<{=�=k>�>O?�? �    N0�0/3   �    �>O?�?   � P   (0�01�12�2�2�3#4�4'5�5.6�677�728�89�9�9f:�:n;�;�;�;<�<�<O=�=*>�>?�? � `   0o0�0f1�1E2t2�2�2�2&3�34o4�4?5�56v6�6V7�7J8�829e9�9�9�9j:�:];�;*<�<=~=�=�=�=?>�>?�? � d   L0�0=1�12�2�2j3�3F4�4&5�5�5�5 666�6�6�6�6�67�7�7�7�7�7�7f89�9�:+;�;"<�<+=�=�=v>�>O?�?   � T   0�0�0r1�1u2p3�3�34z4�4`5�5}67v7�7r89�9):�:;T;Z;�;�;�;[<`<�<y=k>�>�>?�? � X   0(0�0x1�1�12�2�23�3�3)4�45�56v6�6]7�7=8�89�9�9m:�:f;�;F<�<-=�=>v>�>V?�?   � H   /0�01o1�1o2�2�233�3�4*5�56R7�7O8;9�9�:�;k<�<k=?0?<?�?�?�?     X   �0#2444�4N56|6�6�6S7�7�7S8x8�8�8"9�9:(:�:G;l;x;�;#<8<�<@=�= >>>�>�>l?�?    T   t0141@1L162�2�3 444$4;5�5Q6�7�7�7�7�7E9h9t9�9�9:x:8;4<�<=�=*>�>�>m?�?     P   F0�01�12�2�233U3�34�45�56t6�6b7�7�8"9;:�:;�;<�<=�=�=�=>o>�>o?�? 0 @   o0�0F1�1/2�2.3�34�45�56�6�6d7�7K8�8+9�9:{:�:[;�;;<   @ P   *3/3=3�3�3�3�3�4_5�5�5!6H6T677)7�7�7�7{8�8�9l:�:L;�;/<�<=�=�=h>?�?�? P L   d0�0T1�1b2�2r3�3d4�4D5�5$6�67�78�8�8j9�9J:�:*;�;<9=\=h=�=Z>�>R?�? ` L   =0�091�1:2J2M3=4�45�5�5V6�6T7�7;8�89�9�9k:�:K;�;+<�<={=�=[>�>;?�? p L   0�0�0o1�1o2�2e34�45�5�5l6�6K7�7?8�8=9�9+:�:;{;�;[<�<;=�=>�>?? � 4   0�0�0t1�1[2�2?3�3/4�45�56�6 7�7�8;i>n>�> �     m5�5�5 6�6Q7x7�7�7h8�9H? � H   �2!3&373o344f4s4�4�4�4�4k5�5F6l6�6�6?7�7$808�89h9�9�9:\:};#< �    �0 9�9   � D   K4�4k56�6#7�7F8N8�8�8�8�8"9'909r9x9�9�9�9�9�9%:L:P:T:X:\:`: � X   77g7l72:E:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;G;S;r;�;�<.>(?-???�?�?�?�?�? � �   00!0.0_0�0�0�0�0�0222D2g2|2�23@3U3@4�4"5H5M5_5�5�5�5 6s6�6�6�6�677�7�7�7�7�7'8.8~8�8�8�8�8�8P:W:r:�:;R;v;�;�;<@<q<�<X=]=o=�=>>>p>�>�>2?l?�?�?     �   0(0D0J0W0^0c0~0�0�0�0�0�0�0�0�0�0�0"1�1�1,272r2�2�2�2p3�3�3�3�3�3�3�3�34!4?4D4K4�4�4�4�4�4�6�6�6�6	:T:`:�:�:�:�:�:�:�:�:^<j<�<�<�<�<�<===X=d=�=�=�=w>|>�>�>{?    P   b1n1�1�1�1�1�1222V2b2�2�2�2�:D;P;};�;�;�;�;�;�;�;3=?=l=q=v=�=�=�=�=�=   �   )0x0�0�0�0�0�0�011#1�4�4�4�4�4�4�45B5L5�5�5H6M6_6�6�6G7L7Q7X8]8o8�8�8�89�9�9�9�9:|:;;;(<-<?<	='=K=R=v=�=�=�=�=�=�=�=�=>>9>C>H>M>W>\>a>k>p>u>>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>???#?*?/?5?<?A?F?M?R?l?r?y?�?�?�?�?�?�?�?   0 �   �0�0�0�0�0�0�0�0�01113191F1�1�1�1z2�2�2�2�2�2�23�3�3�3�4�4�445=5'656<6F6M6T6`6g6n66�6�6�6�6�6x8}8�8�8�8�8�8�8999 9)959>9_9y9�9�9�9�9;:@:�:�:�:�:;;;;";(;0;6;<;D;U;^;�;�;�;�;�=�>�>�>�?   @ �   00!0-0C0O0X0^0g0s0|0�0�0�0�0161�1�1�1�1�122>2�2�2�2�2a3j3v3�3�3�3�3�3�3�3�3�3�3�3�3�3�34-4�4�4�4�4�45 5*565Q5W5`5q5y5�588=8O8u8�8�8�8�8�9�9�9H:P:Y:i:u:�:�:�:�:�:;!;-;2;b;n;�;�;�;�;D<J<�<�<�<�<=<=B={=�=�=�=�=>>>E>O>[>v>�>�>�>�>�>? P �   �0�0�0�0�0�0111'101@1L1b1n1w1�1�1�12�2�233/3�3�374C4f4�4�4�4�4R5W5\5|5�5�5�5�5�5�5�56z6�6�6�6 7&7o7�7�7818�8�899998:=:O:c:�:�:�:�:�:�:;;1;7;D;�;�;�;<!<N<S<X<h<�<�=�=�=�=�=�>�?�? ` �   000/0U0a0�0�0�0�0�0�1�1�1�1�2�2333<3H3u3z33�3�3�3�3�3}4�5�5�5�5�56q6�6�6�67U7q7�7�7�7-8v8{8y9k:�:�:�:�:�;�;<<�<�<�<�<�<�<===_=>?J?w?|?�?�?�?�?�? p �   0�0	2&2W2t2�2�2�2�2�2%313^3c3h3<4�6�6�6�6W7c7�7�78*8W8\8a889@9V9c9h9�9�9�9�9�9�9�:�:�:;;;J;U;f;w;~;�;�;�;�;�;�;�;�;�;�;�;�;X<]<o<�<�<�<�<�<�<�<@=V=]=e=l=�=�=�=�=�=�=>�>�>�>�>'? � �   �0�0�0�0�0�011@1E1J1b1�1�12	22%272C2p2u2z2�2�2�2 3&3:34474L4Q4Y4n475Q5{5�5
6+6�6�6�6&838K8k8y8�8�8�8<9[9a9r9�9�9�9�9::<:K:^:�:�:
;;;%;-;:;F;�;�;�;I<   � �   �01'1H1j1�1�1�1�122.2X2]2c2�2�2�2�2�2�2�2-3�3�34/4}4�5�5�5�5�566$646}6�6�7�7�7�9�9�:�:�:�:;
;;;;&;-;4;;;C;K;S;_;h;m;s;};�;�;�;�;�;�;�;�;�;�;<�<�<�<�<�<=,=1=6=�>�>'?@?�?�?�? � �   ,0�0�0b1~1�1�1�1�1�1�1�12222}2�2�2�2�2�2�2�2�2�23	332373,4�4�485c5h5m56'6m6�6�7�78p8y8�8�8�8�8�8�8�9�9L:S:L;W;p;�;�;�;�;|<�<�<�<�<�<�<�<=C=b=�=�=�=�=�=�=>>�>??�?�?�?   � �   00>0C0H0o0x0�0�0�0�0a1z1�1�122#2/2j2s2|2�204n4~4�4�4�4�4�4�4�4v5�5�5�5�5�5�566696I6U6�6�6�6�6�6 7&7T7Y7^7�7�7�7�7�7(9-9?9{9�9�9�9�9�9�9:::C:�:�:�:D;|;�;�;�;�;�;�;<�=�=�=�=�=�=X>]>b>i>�>�>?0?<?P?\?w?�?�?�?�?�?�?   � `   00.0:0�0�0�0�0�01111<1=3F3p3u3z3	4'444�4�4�4�5�5�5�6�6�6�6�6�6'89�9�:�;�<w=g>W?   � |   G0'1(5�5�5�5�5�566)626?6�6�6�6C7�7�7�7�788+8Y8�8�8�8�8�8�8�8�8�8$9:':S:c:m:�:�:�:i;�;<d<�<=5=|>�?�?�?�?�?�?�? � T   �0�0<1U1�5�56(6D6`6|6�6�6�67�7�7�7�7�78E8y8�89g:�:O;[;�<8===O=r=�=9>�?   � �   1�2�2�2�2�233?3D3I3�3�3�3�3�3�3�34"4'476C6	7777<7A7�7�788!8�8�8�889=9B9�;�;�;�;�;�;�;�;<?<]<d<h<l<p<t<x<|<�<�<�<�<�<�<B=M=h=o=t=x=|=�=�=�= >>>>>>>>f>l>p>t>x>�?�?�?�?�?     �    00F0�0�0�0�0�01	1F1O1y1~1�12282a2j2�2�2�2�2�2=7L7V7n7u7�7�7�7 88%8M8Z8g8t8�8�8�8�89+9m99�9[:�:�:�:�:�:�:�:;[;�;�<�<�<=L=�=�=�=�=>>>%>.>6>?>E>�>�>�>�>�>�>�>?=?B?�?�?�?�?�?�?�?    000&0�0L1Y1�1�1�1�1�1�1�1�1�122'2�2�2�2�2�23C3�3�3�3�3�3Q4V5d5�5�5�5�5
66!6A6f6o6x6�6�6�6�6�6�6�6�6�6�6�677T7s7�7�7�7�788#8B8U8Z9i9r9�9�9�9�9+:K:S:Y:}:�:�:�:;;/;=;E;k;r;x;�;�;�;�;�;�;�;<I<T<k<v<�<�<='=T=b=q=z=�=�>�>??+?:?C?h?p?�?�?�?�?     0!0'020I0T0c0�0�0�0�0.1`1d1h1l1p1t1x1�1�1�1�1�1�1�1�1�1 2222p2t2x2|2�2�2�2555!5)515N5W5y5�5�5�5�5�5�5�5�5X6i6|6�6�6�6777G7N7T7c7q7y7�7�7�788D8U8p8�8�8�8;99�9�9�9�9�9	;';5;>;�;�;�;�;�;�;<$<7<@<k<~<�<�<�<�<=+=U=]=h=p=x=	?"?0?=?L?U?n?|?�?�?�?�?�?�?�?�? 0 �   L0Z0{0�0�0�0�0�0�0�0�0�01U1�1�1�1�1�1�1y2�2�2�2�2�233)3:3G3O3T3g3t3�3�3�3�344=4J4�4�4�4�4�5�5�5�5�5�5�5666D6u7�7�7�7�7�8W9`9�9�9�9�9�9�9�9�9�9:::::�>�> @ (   �2=3�4A5g5t5�7�8�9;:d;v<)>�>�?   P �   B0�01�6�6�6�6�6
77"7o89+93999S9Z9�9�9�9�9�9�9:: :(:8:A:G:U:b:k:t:�:�:�:�:�:;	;;$;I;�<�<�<�<�<�<=4=}?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   ` �    000`0d0h0l0p0�0�0�0�0�0�0�0�0�0�3�3�3�3�34�4�4�4�4555J5�5�5�56@6G6777 7$7(7,707�7�7�78R8[8l8�8�8�8�8q9�9�9�9�9�9�9:+:g:p:u:�:�:�:�:�:�:�:�:�::;j;s;z;�;�;�;�;�; <$<(<,<0<x<|<�<�<�<�<�<�<�<�=>>>$>>>G>L>}>�>�>�>�>�>�>�?�?�? p <  00%030I0g0u0�0�091F1T1]1�1�12*252>2u2|2�2�2�2�2�2�2�2
33%3?3F3W3i3{3�3�3�3�3�3�3�3>4X4a4r4�4�4�4�455+5b5i5r56@6U6l6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7�7�7�7�7�7�7z9�9�9�9�9�9�9�9�9�9�9::7:�:�:�:�:�:�:�:�:�;�;�;�;<<%<C<O<X<w<~<�<�<�<�<�<�<�<�<�<�<�<\=�=�=�=�=�=�=�=�=�=>�>�> ???"?   � t   m0�2�2�2�2q4y44�4�4�4�455#5(505;5G55�5�5�5�566/6;6C6(797~7�7999b9k9�9�9�9|:�:�:;/;8;A;�;<�?�?�?   � |   0030M0Z0b0�0�0l1�12
3{4�4	5�5666�6�6�67'7f7s7{7�7�7�7�7�7�7�8%9R9`9i9�9f:�:�:�:�:;&;F;f;�;�;�;�;<4<B<f<�<= �    1&7I7�8�?   �     d2=3�3K5�96<�<�=�>?�?�? � �   �1�2W3�3�3�3�3�3�3444+4N4U4�4\7�7(8/8n8u8�8�8�8�9y:�:�:�:�:�:�:6;=;W;^;�;�;�;<$<)<e<l<~<�<�<;=B=�=�=>)>V>�>�>O?X?�?�?�?�?�?�?�?�?   � �   �3�34476C6�6�6�6�6777797_7}7�7�7�7�7�7�7�7�7�7�7�7�7�7b8m8�8�8�8�8�8�8�89 9$9(9,9094989<9�9�9�9�9�9�;�;�;<F=L=Q=h=m==8>=>O>f>m>�>�>�>?(?-???�?�?�?�?�? � �   000 03080?0F0Y0^0f0m0�0�0�0�0�0�0	111>1D1�1�1�122J2O2T2|2�2�2�2�2�2�2�3�3�3�344'4�4�4�4/565=5Z5w5�566F6K6P6j6�6�67�7�7�7�7�7�7�8�8&9-9�9�9�9�9�9�9::2:8:f:o:�:�:�:�:�:�:�:;6;;;@;N;c;w;};�;   � l   X0g0_1h1�2�2f3r3�4=5I5y5~5�566Z6l6�6�6�6�6�6:7F7v7{7�7$8Y8�8�8959:9?9�9�9�:;9<@<=�=H>�>�>+?0?5?   p   0�0�0�0�0�0�0�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6777 7$7(7,7074787<7@7D7H7L7�>??8?A?k?p?u?�?�?    �   0$0*0?0I0c0h0m0w0~0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111o1z1�1�1�1�1�1�1�2�2�2�2�2C3K3�3�3�3�3�3<4D4q4�4�4�4�4�4Q5X5�5�5�5�5�5�5+636�7�7�7�7�788@8�8�8�8�89 9%9�9�9M:U:�:�:�:�:�:�:(;0;�<�<$=)=.=s={=�=�=�=�=�=}>�>�>�>�>???W?_?   t   �0�0�0�0�0&1.1�1�1�1�12	22}2�2+333^3�3�3�3�3�344�5Q6y6�6r7~7�7�7888F:N:�:�:�:;;:;?;D;�=�=�>�>�?�?   0    00z0�0�0�0C1K1�1�1�1�1�1
22C2H2M2A4J4x4}4�4�4�4�4�455+5;5�5�566676C6T6^6n6x6�6�6�677767�7888#8K8Q8l8y8~8�8�8�8�899"9X9]9b9g9�9�9�9�9�9�9�9�9*:;:@:E:J:s:x:}:�:�:;;;S;X;];b;�;�;�;<
<<7<<<A<F<i<r<�<=�=�=>>D>K>U>g>q>�>�>�>??   @   H1M1f13292M2R2W22�2�2�2�2�2�2�2�2B3G3L3�3�3�3�3�3�3�3�3�344 4T4e4j4o4t4�4�4�4�4	5=5B5G5}5�5�5�5�5�5�5�5 66L6Q6V6[6~6�6�607�7�7808A8H8�8�8�8�8�8�889?9z9�9�9�9�9�9�9�9>:D:�<�<=
==)=C=H=M=W=^=c=h=r=y=~=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=O>Z>a>{>�>�>�>�>�?�?�?�?�?   P D   "0+0U0Z0_0�0�0�0�0�0�1�122"2I2U2�2�2�27^7$89/989�9�9�9�9 ` x   �3�3>4q4�4�4�4�4�4�4�4 55X5]5o5�5�5�5�5�566/6o6}6�6�7!8i8�8�:�:�:�:�;<</<y<�<�<�<�<�<�=�=�=�=?"?(?3?9?E?l? p T   0�0�0�0*1/141\4%5�5�5�5q7�7X8�8�8�8�:\;h;�;�;�;�;<"<Y<o<�<�<4=J=|>???? � P   ]0i0n0s0�0�0�0	222�2�2�23[3`3e3�3�3�3444�455;5j5�6%7M7�7+8U8�8�> � $   �0�0�1�1�1�5P6o6�6Q7^7v7�7�7 �    �?�? � d   0U1`1l1w1�1�1�1�1�124%4D4c4�45/5y5�8l9�9�9�9�9H<g<�<�<�<�<=!=@=_=~=�=�=^>l>{>�>�>�>?I? � (   f7�7�899J9O9T9�9;;r<y<g=n=   � `   4282<2@2D2H2L2P2T2X2\2`2d2h2l2p2�2�2�2�2�2 3�56'6	7	=�=�>�>�>�>0?5?:???�?�?�?�?�?�?�?�? � P   �8Q9]9�9�9�9�:�:�:�:�:;;F;K;P;�<�<=="=�=�= >R>�>�>�>�>�>)?2?\?a?f?   � �   �0M1�1�1�1�1�122>2k2p2u2�2�2�2/3;3h3m3r3�3�3�4�4"5'5,5�5�5�5�5�56C6K6�6)717�7�7�7�7�78
8�9�98:=:O:�:�:�:;;;6;N;W;�;�;�;�;)<2<I=U=�=�=�=�=H>M>_>�>�>�>???2?J?S?�?�?�?�?    	 |   00 1D1M1�1�1�1�1�1�1$2)2.2T2�2�2�23_3�3�3�3�3�3{4�455i5s5�5�5�5
6R6�6�6�7�7849>9h9�:�:�:�:
;d;n;�;�;??.?7?D?   	 �   +0N0W0�0�0�0�0�0111&141=1K1Q1Z1h1r1�1�1�1�1�12*2<2�2�2�2�2�2+3�3�3�3�3�3G4y4�4�4�4�4�4�4555>5h5m5r5y7�7�7�7�7�7L8U88�8�8#9,9V9[9`9�9:R:[:�:�:�:9=B=l=q=v=:>b>R?�?  	 �   W1_1�1 2-22272x2�2�23/34393�3�3H4P4�4�4�4�4�4q6z6�6�6�6�6�667?7i7n7s7�7�78A8J8t8y8~8�8�8&9O9X9�9�9�9�9�9�;�;�;�;�;�;<0<5<:<s<{<�<�<�<�<�<:=C=m=r=w=A>M>z>>�> 0	 �   �0�0�0�01)151b1g1l1�1�1�1�1)2.232r2~2�2�2�2�3�3�3�3�3y5�5�5�5�5�57�7�7G8�9�<�<�<�<�<6=>=�=�=�=�=�=I>Q>�>�>? ?M?R?W?   @	 �   �0�0111O1[1�1�1�1�3�3b4n4�4�4�4�4�45 5%5N5�5�5�5�56 6%6c6k6�7�7�7�7�728>8k8p8u8�8�8�8q9�9�9>:J:w:|:�:�:�:[<�<�=�=�=�=�=�=�= >%>*>e>m>�>�>�>�>�>.?7?a?f?k?   P	 �   >0J0w0|0�0�2�2
33393E3r3w3|3�3�344=4B4G4�4�4�4�4�4�5�5666�78)8Y8^8c8�8�8�8�8�8�9�9�9�:�:�;�;�<�<�=>?�?�?�?�?�? `	 p   �0W1^1�1�1�1�1D7H7L7P7T7X7\7`7d7h7l7p7t7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888o>{>�>�>�>�>�>???   p	 d   ?1K1x1}1�1 2R2�2�2b3w3�3�344474L4�45H5�5�5�67777R7m7�7:4:�;�;�;�;�;�;�=�=^>l>�>�>?,? �	 \   2�3�3�3�3�36;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;p?�?   �	 D   �0�0$1)1.131d1�1�3�34^4�4Q6�9�9�9N:<<\<�<�=�=>3><>d>�>R? �	    &1D1�4�4*9N9�9X=]=o= �	     (0-0?0�3�3�3�6�67H8M8_8 �	 T   80=0O0�0�0�0x1}1�122/2�3�34�4Y688h8w8�8�8�8�8�8Q9Z9�9�9�9�>�>G?]?�?�?�? �	 T   00050:0�0�0�0�0�0G6]6�9�:�:;;;�;�;�;<J<V<�<�<�<�<�<===b>�>�?�?�?�?�? �	 �   �0�0�0�0�041�1�1222�2�2�3	494>4C445@5p5u5z5�6�67"7'78$8T8Y8^8"9)9�:�:7;C;s;x;};G<S<�<�<�<�=�=�=�=�=�>�>�>�>�>�?�?   �	 �   000�0�0111�1�2�2333�3�3444�4	5�5�5666�6�677!7�7�7�7�78�8�8*9/949�9�9-:2:7:�:�;�;�;�;�;<"<�<�<�<�<%=,=�>�>�>�>�>�?�?�?�?�?  
 l   �0�0111�1�1$2)2.23'3W3\3a3+474g4l4q4D5P5�5�5�5T6`6�6�6�6{7�7�7�7�7�8�8�8�8�8�9�9�9�9�9�:�:�:�:�: 
 t   J0V0�0�0�0>1z2�2�2�2�2 3$3(3,3034383<3@3D3H3L3P3T3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3$4(4,4044484<4@4    
 `   5�5�5�5�5�5V6h6�6�677>7C7H7�7�7�7�7�7t8�8�892979<9�9�9:4:9:>:�:�:�;<8=?=>�>G?�?�? 0
 l   *0/0401�1�1�1�1�1�1�7�7�7�7�7084888<8@8D8H8L8P8T8X8\8`8d8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8   @
 �   H0M0_0�0�0�0E1�1�1�1�1%2+242I2�2�3�3�344"484�4�4�45(545@5V5�56&6^6c6h6�6�6�6�6�6�67�7�7�788�8�8�8�89K9i9H:M:_:�:�:;;�;�;�;�;�;x<�<�<�<M=V=!>�>�?�?�?   P
 �   00.0D0m0z0�0�081=1O1x3}3�3�3�3�3434O4y4�4�4�5�566-676V6�6C7O7�7�7�70898c8h8m8R9�9�9�9:@:l:�:�:;;#;e;q;�;�;�;Q<�<�<�<===d=�=�=?? `
 x   A0H0%1�1q2!3-3]3b3g3C4�4�4�4�4*515�:�:;	;;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$< p
 P   �5�6�6�6�6�67)7Y7^7c7�8�8::>:C:H:�:�:&;+;0;~;T<[<m=y=�=�=�=�>�>�>�>�> �
 �   S0_0�0�0�0�1�1�1�1�1�2�244�4�4�4�4�4�5�5�5�5�5A7M7}7�7�7S8_8�8�8�89@:L:|:�:�:R;^;�;�;�;<�<x=�=�=�=�=�>�>�>�>�>k?w?�?�?�? �
 �   �0�0�0�0�0�1�1�1�1�1�2K3W3�3�3�3�3�3]4d4�4�4�4�4[6g6�6�6�6m7y7�7�7�7�8�8�8�8�8�9�9�9�9�9�:�:;;;�;�;%<*</<==>=C=H=> >P>U>Z>;?G?w?|?�?   �
 �   M0Y0�0�0�0c1o1�1�1�1u2�2�2�2�288B8G8L8�8::N:S:X:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;   �
 (   (;-;?;e;n;�;�;�;i<�<�<4=@=>>   �
 �   W0`0�0�0�0�0�0�011�2�23+30353^3g3�3�3�3Q4Z4�4�4�4�4�4�4�4575@5j5o5t5�67$7Q7V7[7�7�7�7�7�7�7�7)8.838�9�9�9n:�:�:�;�;�<j=�=�=:>^>�>
?.?�?�?�?�?�?�?�? �
 �   000L0U00�0�0r1{1�1�1�1�2�2�2�2	33<3A3F3l3�3�3�3�3�3�34!4Z4c4�5�5�5�5�566;6@6E6�:�:<<�<�<�>�>�>�>??R?W?\?�?�?�?�?�?�? �
 �   0Q0Z0P1g1�1�1�1<2E2�6�6�6�6�6�6�6�6�677777 7&7,72787>7D7J7P7V7\7b7h7n7t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78
8888"8(8.848:8@8F8L8R8X8^8d8j8p8v8|8�8�8�8�8�8�8�8�8J>a>i>�>�>�>?J?   �
    �?�?�?       _0   0 �   1114 4$4(487<7D8x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�> @ <   �0�0$1(1�1�1�1�1�1�1�1�1�2�2�2�6�6�6�6�6�6(;,;0;4;8; P    044484<4@4   `     >$> p 4   \9d9l9t9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9: �    �1�1�1x8|8�8 � �   (1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�6�6�6�6�6�6�6�6�6�6�6�6 77777 7   � ,   x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:   � �   �<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>�>�>�>P?X?`?h?p?x?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?         082L2P2T2    l   @4D4H4h4l4p4x4|4�4�4�4�4,>0>D>L>P>T>X>`>x>�>�>�>�>�>�>�>�>�>???(?@?H?\?`?t?x?�?�?�?�?�?�?�?�?�?     ,   000 0(0@0L0d0|0�0�0�0�0�0�0�0�0�011 1(101H1`1d1x1�1�1�1�1�1�1�1�1�1�12 282@2T2X2l2p2�2�2�2�2�2�2�2�2�2�2�23$3(3<3D3H3L3T3l3�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 99999999 9$9(9,9094989<9@9D9H9x;�;�;�;�;�;�;�;<8<X<x<�<�<�<�<�<=8=X=x=�=�=�=�=>8>X>x>�>�>�>�>?$?0?h?�?�?�?�?�?   0 �   004080T0X0x0�0�0�0�01181D1h1�1�1�1�1�1�1 2(2H2h2�2�2�2�2�2�2�2�2�2�2333@3H3L3l3p3�3�3�3�3�3�3�3�344,404D4h4t4|4�4�4�4�455@5`5�5�5�5�5�5606P6p6�6 @ 4  0 0<0X0�0�0�0101p1�1�1�1�1�1�1�1�1�1�1`2d2�6�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�:�:�:�:�:;;;;;L;P;T;�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?8?<?�?�?   P    �2�2h6�6�6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          